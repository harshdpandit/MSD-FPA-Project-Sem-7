PK   �fWV9!M�  A    cirkitFile.json�]]�㶒�+Ϋe�"�yۻ���	n.�3C�c{�Y�;��`��%�-K�TRU�d����m��yx��,�_6�����O�r�[y~<���7"�n>���s��6�n>���i��9��a���\��TٹL��m�y)3��e ��΢<�cSi�*�EiX$�>܇�7o��秏�N��x٧�
�X����H� љ@XVd��{�l���2�eTU�@�Fi&�@�2�*a+-ӽ�]�� �G�.b�۠!�]�Y�d���0�T&+B���ľ���f�Gu�Q	J�y`�,t�� )Uh��DU�{�i,3x��̂�*�@��bc� ����R�����0��ഡ�J�����`�2��8����T	�^�u�J�T�B�K�T	�ޒu�J�1Y��p��u�J/���*�``h:E:G�E�t�$� -�IZ�)�,����@�b�Mqݜ�@輿�6�/��͕��A�.!���]ؼ��͉��ȅ���ma�aZ���IYڞ��/m�'����������,�l,�kA�z��l
�׌��<q�H⚑�5#�kF	[[�+�����SD�)��Ağ��"9h*�t�I]Q���/�J�:�D:��w�An�M3��B���`�^��Z�z��}LoJQ&Y^Zk�Ԫ ��	T�L^(�r���3�z~�gF6�9U�G&h�/$�)!h��ha�Q7Mt�� 1"l���\G����/�C�RNf��/��>�G��z��Zͧ��|�gA4�rY��V����띠{BR}�Q´�r�0�uL{"�'��<C�9�9$�z�z�R�\F`J���iZe������2��~���=��`1�'��i>WL�	�b��vbP��2�܎i>����(
q�U��V��ڿXp�Ӛ���������� ��!H�J#��_,���łj�_,X��M�o�u��3�$�v>P=��2��e����b�T"������0d��4�~�w&B���b�	]��r��P��q��]�Z��RV����LOY�|d�lI�KA���滰�GӈIP�*��Q-Ȥ�49M#ť��:+�G#&Au��FL���	����<1	�3<x4bT'��h�$��Ca�H&IMn�Nl�-؈�KR��äw6����
1���߂��}���_���)t��i��D�*TF��A��LI)<3���'�x�؊dJ1<����K1< �1ߊ�Kڅ2)(bZ�UBb+�d<^]���A�L̃bɃbɃbɃb�CĒ��%�%+++&W�ŪFqT�����Q��8O*��Yc�A�Cc	Rj�$%X� c��u��N�Md�"��6RJ���|Cl
ܜ���9��"�R� �b� ap	gRZ[���9����L2m� ��!�� S�8��B�86���I`34�L�d^��y�!�������� �E]T)�k�i\��'2��u�	��5�6[�A����n1H�]�L.)�K ��Š����jq�nv	`����Dl&��#a�����4����R��D�	GO$�6�I@�A16�gz��s;Lyαy����!��X>]��=ǆAPs�â�����E#&A�Q�FL��c-��5Gd,1	j��X4b�ݱh�$�9dшIPs�Ȣ���x��"�X����x[�7����G'6�l��%�=�щ����$�ȱ�K�96t)L�ȱ�K��fE�]�Ǿ�ȱ�K�ر596bx��#�596bx �c�596bx0,x@,xP,yP,�8�ŒŒŒŒŒŒŒŊŊŊɕ�A��A��A��A��E1:ǆ.e5����96t)<� 2ǆ.���96t)���̱�KAd���˃^�_�ͱa�`�_�ͱ��α�K��nl�]
�.�����Х���cC�2O����y����0�n�����%�α�K�]����%�α�K�]����%�ϱ��α�K�/:�fR
:ǆ.e���96t)<�2���96t)�E�u�~i�b�?�o���|>������4/���?���y��niJ��~Ky�4%b��Ly��<3��֔w<S"xJϔ,~�m��H����}?���%�O��{K�K���	'v��q��W=��DVB�i
����� �*�,7��2�l���ۻ�Q���|ՠ�M9�G���{-
�If����'���-4����?�Ly�=i7�2��s��c9�yR��SkR���ѐ�5HOM
s߿�FI����7��c11��Y���uNR�=� Q/6�XjR����
��)x� �� 9Κ���[#J�z�ůê��%�b1(&��!�h�#�Z�o;�3��Qb$^�(|S,��9b~1H���Ü�1<�z�Cyj F�/IO����PS�{:�a>�7G��ƀ�Oj�*�?�� �& ����������SվM�����P0�� ����^0���~ݞ�YDs?�����)��J�E4��Z�E4��Z�E4��Z�E4��Z�E4�%�Z�E4�-�Z�E��5�,F�������@���O�2��T=8T0�(]F{番�
"�X�M��%Q�������]�[(�P��=uvna��mZ�~`U��i`�
�rH�K�s� *�\�<d�*�����t�[����Lf"��,F��$�(��
[I����VR�SR�SR�)���HTT$*�I�"���ߣ/үODC��)�8U8E_��=-{e �����}��"?���(G@#�q�SΡ{����=q�_��#�}J�Is���Oi?��P~ze���^��ThҔ`���L:5�{�$ E���-a��~$�`o���{���~
aػ���S���ߧ�Fz��}����#b����_-��}�w�)�'����Oi?o��|J{<����)�L�}%�'<�ѷ�q��z�����qO���/ͷ�����GK0b}ؑ��lѡo���yBf�u���y�.����v�]�s(\2
�t�(��|����ͧ����M��� �	�s���Q�'�~�Q����p���^�=	נNg����e�ҵ���t-�k!]�ZH�B�ʵP�:�E��T�t)�B�����??4�D�w0�.��A�g�^I��PI�����R1lx�*��Y�FQ��nU�a�%�Ԭ�cyqc�`��91�7D(�Z�]��ʃ�v�(�]���y�U�ԛo{��L��/R`B��#�Q2�3D�����x����W�U���ʚ��/�1�<U�,�º�+�C�է�kܒ��m���el�w���6�s�~*RƆ�v���{e�C���]����Q^��p�D�EbX$�"9,Rm��H���(����l[d�Eq[���(��h��p��p�C\���qO��=�����xqh��H*-��H%�oa�aUe�B]Vq�%�)�����J���?���ı��&K�=x��>���'M�BD�7`>~�^\�����Sy�J;���<=.��*RʝN:���R;+�DG�x�`�
�\W��V&�T��*�m���U�q\��B�~I�y��o7��4O�6�q>��}��`�.ښ(|��}PQ烼��=�ݚ�S-J:��u�&�"ӭ��T�DtK�N��;%�vK�n���n���dw>��^m��d�{��`�47R }-BO�v<G
��v�Z���i�4��&P��j�۩)���ё�IVH$R^�����$��W�.?_�������,k�;G�#Ĵ������j>^·�@�����J���҇'�����t< mn����?�dn�T���<�rx<d��s��O�s	�tB*����4�<��+o��w�=k�/EZ�����p,�\x�V��"��h)�J�k�H����Y���*� ��E��$.� ρr���U�����gd01}>�(o�s o�Va��k�G��X`Ă�4f��v)R��B� B˛qk��a��j���?~�4�o������Sv��#!��$2Qܮ�P�ߡw��m7��.&lQ��+�i
1J��S*� 4,�oY%C�qJ�����뇡�f 	]]mU�HC�@�Jq��%vJ�pӀF �T���&6lD5N�X�(��H-DWv�^lv2N�N��9Skt,�V!�P���&a�0�Z&�9e�U��Z��W�\��L��zv��ZҘV��jX�PK&���r�\�kS	c	�\h+���^�?2j�����P��H]�)E����Z�T���X=��wM�gy�����Z<��s���Gf�t����� �����6�/�8�[��N�ZD�Ś�2NY�
�2m�@��
X� �UV�63*����:#�1N�ob��ɭ2�(n]T[�������
 o8������6��N)mM����UԱ�ed�6Y !O�4����J+��0�j`�Q��Q)N��-���xQ-��-�'�j]�6q+���I�UP2�����6q���Qm������Tmc�w�I�Z�P$��ĉىDذ����(eU����]�E[���^�lc���PQ3�#��Ovk��^����!�����*gc�FFm�9p<�;b�e�B@D�
�)�ȈPF7���7h<h��F�r�IPD8����^>�;@Wq� ��8�$���M�"�*=�u
�PJA_�z�T�F�`�7����IbW,���Vn�����T �gga�e4[�ܽ�L���}�T����DQ ��C%x�idR�e�d�ԯ���*�"Z���V5�TÝ��2��6���a���Ûh���V���L�������@�P ,�*x�:�A�*�����׵5�x��ev�de��PvKT��i<�Dc��mX���E�]N�Fl`t�>���ں�����Æχ���I�L���n��T�o�8C�����m�������CY���g�ӹ�\���P~�O�c�q��ݦ��w�7�6�;�ƾ�l߁㔞/?�?u���ZXy,&E�rbjQ���Ϝ��������p���^>Բ��{�n�(~�~r?������[�߻0n��������	�T[����ZI���_�m�����(�`�l�a�@5,h����4�h|2U�kd-i�x�uD0/�X�U�~�I�=��&qin�܄�������87�*�mb�XgX�a�q	�|���-P��uV�>�����'3��ky��`(e��U�<H���G��#��Y�x��<�%�<I;:�@SP�z�Y�~���mk:
Gk�#�\Y,��ri�������̨UȨ7�W�o��ՒQ'$�ry���/��VhE*8C�D�9=�<>e|�Vs	��.��Vw��G;����[�D��N��jB�pP-��i�ha1`�U�bъZ���g�͔�Ĕ���Z��6
K�,������{���=�%�a(c�~�}��i־{���d�αؽ}��sX��� ��.�On.�\�N��`1(�c	$�f�'�K�ٽ��X�,Pu�3�PЫf�f:����.����Aӟ�Zp+_�Y,T]L,1
,�j��䰚��Zr|�>���lʅQ�NW��y2�ّ1X -�n1���A�N*�=��6U�9Ũ�ƻ>��|аEq��h>��}��Zh�8h��=�Rz�'S���j��N����r�Ť�49���|�r/�K<��J������Yͷ+'��]�o��^,���J���m<(�W��pM5�G15�p�Fɬ�)j��aZ�7}�����2�=`X��6�3��}�� �_�x���d��xp}w䀭ս��\�{se��8�r�I�D�-|�R͆v�t�2�jU8ק5�����մ� �wh5��㟸J���ҷ�0pZft,��zDt��Ӟ,���-�w���ƑUi���	�F����@o.Q���GM=B@V��<�@��TU(����7l�,Ѝ�7V9�t�ځdE��.q����'�OQ�|���gXKgbU�����<����FgxO�LVT�l�5�B��Vk0���~���^��!}xܼq�{�?��,���҇��>�p)?>��y�u��PK   �eWK��"� I� /   images/4354f621-4db0-4aaf-904c-1fa28584b36b.jpg�XSM�/�C�R�*H���4�*�H�JB��������һ�t!6���{�"% �	`y�������y�a��=�Y�ff�̚�l��M�!�
���x���a�    �	�'��� (HLH���t1�( jR�A�M�$Q��t�ݑ!_�v09?7�jO�.��H���(S�T)\#]r$�N
9H�l�e|.Sn�#��ȕm<I	 ��v�O��Dl���,Tddt��� �(�+��@��̽�(d�72@@GG@����ddU�de�dd��T�d�H����OR��&�^��f��A�d���[nGW2�AP����e�7��IO*�r a��m��	�[y�H|���z���;�c$L��?A�4	��R�.��B�cGƂ$�@В"$|#�bk��U��8�<��YVF��w{)m��))�����$��d�^wf���$���w��ҷ1�(���S�!#�N�˒0#)"�)�N��'�tSH߶�TV$�=$��r;9o$�^w�c.���L��zw;�+�NN�W_�C�_�]"����]��i ���QT��#ِ���ܯ�������%-eU$��<��%��-,�L ɫ(�(ˑ-D��Ck��BB�m�wa�-y�n5 �Y{���������ɂ���bۦH|�L��.��N-?Cbq`�Zf\tL q`ڊg�"�~�"�@KKKG�@G����~�>f�}�ll���8Y�h'�{1��������������N�1�oga��@|	����G`� @�
�����~�'�AHZR��h�������������D� �&�  J��������
� OJdS�+K�}ҍM0�5����Ǆ��Y�r�W:ߪC#�`�mt�����!�[Vz��PJ�۬?þ?���=��/z;���;o;Ɨ3J�:���x�D'f��w}]U6��
���U��=�c%�I[�-�h���T8(����A� �ܹ��d^Y�~�v:��c���(BMV����6�i�=���P�ϿT��5���` o��
@��Cq����hd���	�x�Q��@�8w޹�A�9t\F����:>��rr�|#܇���:7�4������b��ax*��G��g��:F�����y�̄�?� \V�i��
v�Lg3�J�����&`��$����mUV�w��t��<3���	��Ws������)$2����ܜ�Y�/[�V�� d~���\3�*1py�`.�2�fc��H��ȣ΀a�x� Raڐ�x��J��i[����a.��nb&�s1"��S��B�x\�5�N��f��;5)��*�N�E_�҂/��]�ޥޞYӼ�ΛDY>
q�it
d<�4�H5�Ux҉��ƨ�IT�C ��O9̙$"���u"zz�^��1���H��(u�g0���y`��YOQā��u��C��C��D���kp�hV�3[ov��I�w>p�����oz&�[�2YZU2S�j��I4k�v�p��O)��O�Ƒ�����W�}�~1�4����7S��4��Q��^XIQ�K����4h�w�<�͵�Zeַ�bO�G]�%TS]%��4�����ی$��]����#3� F��EeE����|��G��D]/�,�ȟ�Bx� �Y�p�Om��H��^��y�G��(ҦON23oz�3�v�9��k+������k.��l�&�o�������z�?L@�N��DEt���G)��}��#�)؏94+���g��И%`6����N�z,Ϟ�z���*��}�u�h���n2- ��u��<���ԧ,AҊ���$��R�d�nv}�����/��x�Xr�tW��\Ȩ}�z�,լ����t�a�^��J2��^�y�j��]����6lR�)!ѻF���'��شފsJ�έ����p����LI�����ǻ�M'z�媱zS�"���L�>J��$�!F��+y�Q��WjlzK���]�ׂ��7��@Ҿ���S��L����^�H�(/���|S�śW���R���F=%�����L���V�k��˸�sj_��VkdF��.{lGV��d$d����-H�n�iK�&��W�"/u�&Vtԏ��C��.�$C�v��L����j���[�ejA ӛJ�C�;Ц��E.SD���W�k�{��o&7�6�k��혷�Ϳvr���,ڕ�8z}e��h��R��ʻ�
�[1�����/�"N'���l]ŧ^W���g	{�ŉ@+f����IZ�����v����e{�|����JTim֔��4F��R�|���^K��e��yP/'�@�l_�fu�A���e.^Kb�Z���:���T�T��Ä��`[������%�
�I��WM��1�����"�$��I���"�T���HcӼ+:�_��vÐ�oBã��s�!�ef���+�_���\�����۔��a1X��N&_�����p(�YP��wk�ш��eG��P�� ��^�V���ۃ�x�LN���v��lN��+��ӑD��O&����O�-h-�ߧ�)}�ؿT�,�����X��� ��Z4��땽�s/i��V��X�}�Z��Q�¼9��W���Ww9��L�Z��Gڜ���B_�@:�G%M���OA�z��?�%���.���nֲ
���>��4%ޫO��Z�M�s��t�d��F�S1����i~��(3������D�˔���sw��� ���s�]�+�Ŋ���.i�!]1�UV�r����Q��v%���b���K��6��c��ܾN�'��Z��Z�������Ծ���M�]��*������ՙ��cgc]&U+:mV+��%�K�Kr�:�>�$�/xM�l���,�����a����wxu,Uc�/8��v���}͖�U{��R�YB�H�M��N��fO��]Z�1����ȅ��-����
��KE�u�.��&�iD�`��T�(��X¬������kU'�rGYBR�+�Y��-�{�5�-�oJގ�I��d�v��.,�+��?l֛�����F�6����������7�'�}]�b���6Or1�~�jܱw�)��+����E>y��N�%�܋+'��u��}�C�����&��S]�q��u��K.�dȍ9�/��<]���+��4�m�ݸ!!*R�B#*�y݄�\p�z��5Y�k��������iB-�7���ɗo��J�.w�Y�q���:�7YJذI5C���%���AQ�G+)5��S=��N[F����z2-VZT�1�8�w�<#|�@��Vރ�\���]���(��.O�L�K���u��2�2���0��]��|{�<��ޚ�2x�[��ZU��=����6�&7�\�F��G�/k;�]�A��W8���0q�xF`[�gg���8Ty�Z��TN/-
�	X��V�ZNb7EK�=�􏽬�os�r����@7�yr��P��_y&�~�껑��l3��!ھ�͔T�6��*�P�������n�wQO�+�r�}�-]�(d��C8,����r3a��:�Q������5�_�JrVF &���W4����Y2�%������
O�%�:�R%-�t�=캕���w|kt��2���E����o�tg/< f���^/ +�56�Z��U����Eq���؄�B{�����稸���j߄����K=��oB�7�rZ�&dh{�[�NO�G��g&�4ϯ�d��bϾ�q��t�)g�i�S�xT<�CA���eս�e5q��p������UQ&�(�WV�G�9�1�s�^x��eJ��W�I�n�st�v�#>����U���O2+&􂟭��_��;ވ��ɖ��y�J�L��O���~�kغ�+=�<:�&��k��|���̴A_�y�A��%��ꋻO�VpȒzՏ�����>8�c�³����=�ry�m�Ȱ��CI��QZ���C��mR��ۮ���u/�݄�zM���\����:�?�-�:���E��E@0Ю���;+�gN4V���p)*�p��3�<��0��{vEA5Ϗ��t�Z�/���M�jYiꨄƖ��<�e�-�l��Xf���9��>�9W�(ΰ#�j�Jt�m��H�̶U�����͈ˑ��hN*�W%4�*�����qغ��<؄��]Rfޥ���Ǵԟ����S�>��_2'�bD����B��x�2�F&`�� ��W��X��q����F��v�6��N���(c�Kf|����D�ߗ�Y��]��fj�l��o��7[��k�Q2�JT]�g��iZ�8衍��q�]�b����6�~�����%�?����/���GlBL��HK��R]�V�����N���l�Y����H�$��}���֘�>��|���[\~��U��F���|ة32mY2����k��&'/�qWq3M�%� ����n��J�L�=���t��aEm��qh\�Ca/�Ji_�k�i(����L�v]'����MGI<���yB�������4�jV��m�a����S���2�n���X��j=�U|���tB�z��%�B�v_k~���1�9�@�
�2�M\�C�9��f$��4qas���|Q�,�B�6k��i�zq���gs-y=�FdM˦W��q�>��I�w*Y�vM���`B+��+��PeWyH������ދ�F<z�g�0����_Fyn�-n�,�{m���q9���5������el�{���o��
j�c�E�#��e����V������(�5Lf�=di��1�?^�|� t)�F8�n�mg���ۊ�6C�W� �Y�e��=Q7�6
S�6}���5��O�{z�<-w�ݠ���H5���K��ڦ\�xCu>���> k?��#X�7���i�v�n|�ehԭe+�O�Ճ�7�N�������}�5D���{����#�#�-�]L�^#��:�F��`..�h�)� g�l��0�𐎷� �3Nvo��_f'&�O?\���)��������JH�vysI���1k˷��M9L���ﬗ}<Ҫ0�}���O���پY�گ������n��~����/K~c(W��W�6�r��~4Qm�N}S�ֻOi�~E��Nl�,1��]�׌�S�.��X��y߭�P���_~��<*e�m_S�؇�#�*�eyOˠh�dZ�U74�f��zTs���)5��]D�s�~�)��<�S�K?jƛO%���\~`��\_��yOV٥4F�ߙ��%ʬu�?��'tG�Yo`�0�^�\8fE��b��5�0���%6����A�D�!�^E��u�R�׾���[�c�&6x�����~ҞRl�II���<r8�&��者�ȍ��u��]���Z���w'�V��s�*%Z*�(Gq=.~	nC��_��_|C��"�ü�
�Ϟ��D�N���g,�0���OU��J>a�*�H3�y��N:ߟ��O�K��Y��E>��q����Y�ױ�Ւ�D����e���Ь�?�{������3�.SIs�P�/J�tBl"i�~_/H>͏��c��@�&���J���4�d�:c�!42�=5���ô�buJY�@7�93ҥo"]ΰ{��l��2?��̙�U�ŧ��D`��*��FvA�{7CL5��ZOK�e����1�|[���{�ߔ*G7B�"ˢ��lh�T��~s[;,u���pLA��ڛxv����/�D`/#�G���lhϻWh�)ƈ2ۄ.�^��n8fb�W,�P<5���SR�}�k,�?��P8�"�i�]������X�]��5]��n)Zo��.� �R�>���o��
.�n*��vm�Ma�?k8�!�y��+ز�WE��i>\�BbE�	
�<���πi�]����Ux�4a�2��I��:6p8��\m�4Ψ���2l�r������R�Ů�o��f��͈OIWYy� eں�P�3�뱷9��z@������|_>"`��׀�<�q5;ϿV�q߱�۵���I2�w4��a��CjY��Z&�fL�ٌ���jj\ulHn(�-k^"	�`F�0K���"�"�l|#��E��u���d��Įߖ�����u@ư���Y�����_�JjSb��!Vx����f�q��̢{�W�F���s�ϐ�J6���W�������WR����5��G[p\�+c����F��됛��S�� `�'�s�ך�зn^;��iǚD��!���_�?M��?q��Vf�Jņ.��#��f��r/�gMi)��=_/r�~s^���"�ʱ�P$�iu���7F3��@j��� �_�iug�V�`e� ���4�
j��j0|Z��C%#�����%���<QF��Қ��Nh�I�T#K�����#�=\�dR�ܯw����6*9L�}��j���u�F��6�B��7��"�ܠ~���n�#g�h���Oa'�Юz��d�'|�-8�;᫛Eȿ�i�j�I�����[�u8�ei]<��5/�l��Ј{sM����t��1OH��Ӟ�5�?/�|�#m���͌P*�Ö�ЈM!�;q�`�����|xcߙ�r�kY�yG������~�w����|�ų9�R~�I��]��3����;+�/E�|l��lUC'��}A�9ݽ�W�2"����y��qڽ�N���Hʺ�Y���c	�؊&�~���bn%�PVC��������v�TS2����)��!�c�xIA}V�'���p���}�"-r����C��_`Ib�%�q$����7N�$v�ađp"P�lNZ� +ڰѱ�;I����h�t��)" G�H �3�'��36����I���Q�o�m�L��xN��[f>�������9��Q�[7�p���x3���l42�'nzf}�%��S���s�ެ�w����94�}5��o�aF>�S��j=�b��=�"��z߻���2�
��T�6��ok�a*���h��P+���Ѣ���	[g��w3�;`��*���8�����D 1�^.� e��qB]�S�������=�Nw�Z�7&8l�t|���]_x���{k�����D��u8#gy���'V��*����6}s��5)re�s�˘�p�b�dd�.V*�>�!O��4�Ըd��nꮩ����ܵ�]5,Uz}�5��������wЎ�6�b��P+�<����=�])�%�A�YY���:xy(ռ�:h��}yG=��@&;�u��[���>O(�{j8���8/�����u����di��)�!���H���G����%>⅏N1  ���k1�Y�\L�M�Pu���\s��Hs����z]<10^	Y�"���J��\F�b���{��\3*�S{qAo�w~	)�i)Ҁ0������S��a����H�&���i��ɢ��� �`iJĆ��-��#W Sx��չ_]�d�̻U����U?�{(/Ğ�f1���_��iP�&���W�|�tD1)���@��/j"�C���eny�o��S,P0��Ro2��Sl�`R�-��e�9�6�*��ʳ��A��fL!�i�R6i��>��=8u9�૵CiK�S�4�C��y�x���J����������h�LO0� M��?_D�D����U]xէo�����S	D-+*�C�;�ϲ�z?中?�DVQ`5i�S��j�P�.xh���U�ip�y|�Y�(��"f.3n��. ��`&"h8Ɲr�r����h���%�c�K������y���O���N�<,v�i*n�0e0`�_����]xFn�ܘe��$���/�>'������	��QY���]���H<����㌳�+)��5u���{�qLl-i�9�8K����	6��%�	�;��h6F�Z7ۊ*>�.��%C�k�ǈ6C#"pzx��b(�E�Xc�W�]ք��D����8,8�4������@SO{%5�v�")j��x�0u�A���O�)8Y��۽���w_qY��BZ�$�H+XSp�͎t��r���3e�����h'�؝V:3p\ �m>����6�`���C���^✨�o�y)@嘡	��/� ��
) ��=��B�%����(�R��BeY9	���"[�Y"�N��2~��e������4���n`��c��잀 ��
@��m�<e�D�mI"P0��o��^��y+��OY����w�� S7����կʶ3�!���0:���J�����rl-�%D�+�g�c~(Ď�h?�b����������v����)$��ƽ��, �D����I:(�O�?��_�`��)A���w���/�W���+����+B��E�½v���j������Xxx ��Zȑ�~�A��x���]�X���5�/d���c~Ƿ�Cm�����,~��C`P2H����̽̃��:[� �D�]�V$��;�%�o�oղ��f�!l�a��%����g�1�,H:C�PH?$�k'���
��-|���L��3���/6�r�s�:�gP�����V��@������a @ܢm.%��<�lŹ�/m��~���%ʲS�/'�-ٕ-|���$�����;��9����őۺ; �/���]�7g��[8���J�Ir���i[}A���[�O��}���O�qn2���~;������	` ��Z�ȓ��ޱ
�7y�#�_�{� h?���{�ݑh�G��^(J���d���܀�K��/��V��ynũ��|��`?c�����4`�!�f+b��G�4^AHt�_X�� /�_k��%9���gtC��0,���:�:�s���&s�);K������������{��g���e���F�C�21�����d�E������������'�ܻ0O7��:FB����O�_���{� ��At.�v�c��j�"�� �X���8z?RG���}kA�7�� ��/�%���lΐo�o>�$!�V�,���G�h !A>�	�v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v��v���O�_�zK|p뽨%��(�%)3�x H���9�M�(�����\{�	@�~z�Pn{}�l}��Tq����
P��FK���5KA���anҲR2��QHX�C	�ü|��XAA[E� ����� �e��4U��h
S���������ja�[���0�--(�%��kn���\@P�R����*(�J�*�*���������������S�QU�U�!ARmA�j��;u�b�;�
�
��ByI˪��J��I��I�$$�O#Pna��`��%��A>[�l丛;������_��m_����@�mU������aT0IV��l�Oſ/�W�_* ibb�����K:���ϥ�����`$:
�!�)D��f����<�놂i��$%ee%e�~~�KBFEMFf[T'�BY!�~?���?���8��K����N�$S�pC���
x@�<�A�n�����y��}`^�ǂ�
�m���ZC*F�O����y��Ǐ�lapL�POGIVUIIRNJ�OA�
�:{��
���"�Qn�#�� �#���&sS��S������K�++�J��*�J*y�z()�@a��*?��"�h����������\y�n�t�'�4��wf�%,p��lٔ��<WH����a���ۿ�?���O�z[,�
u�i{���_��v��<z҂Ҥ�H�n���6X�_փ�,�"�%�su�إ]ڥ]ڥ]ڥ�����A�Z���~���H�Js3}Cc��9���>$ �#PA�}���� �'���Y p��X�[m�����7��_h�k۹�]򸹀 �F�Ѐ �Ϝ��=H;�H�~�� 2����'c
��2{IA�$c�m|dKfk���?��:x�{��[��&;���I8:�J��O���}H�|V��� [^��(ԛ���e�� =�R Z�?���:���8��-  =�����P(IsҠ�y�)���`��[���6�t����$��n���۟A�h���;9� PY!�͍�<�� P~	 8�~� 3i�ʚ�h�^�x���A�����K���Q���_�#���/@�7(�1$L�0�5��qƿ���#=lؐ���En������?��a��m�&[:`w�X���\@ɶ �zHJ�7c:�<�l�'��~���E<��u4б����B�ӶN�P� 3�p !@�� e@���`�� ���  8���X�p���@P� ���P| Z�N�� 3�7`X�@4 F��I��@* M��d����@ttJ �=倊A��W�w�VP/h4��S�)(�)�(QHS�PhSQXQ8QxQR�S\���H�xB�OQF��E'���
 �s��%�*`���	G�c���'�Bp��ς�(�)�((%)�)�SZSB))�(�Qޣ̦,�|K�N9J���@�H�K%A�FeHeG�EJM�H�IUJUG�I��j�����Z�Z��8�=�/u�5��E�/�[�ǨWhhh�h$h4h�h�hP4�4wi�i�4m4_h~��姕�էu�EО�M�ͥ��m���]�c��S�3��;MO�NWE�L��n���^�^�ފޗ�}2}!}� �Ҟ={���9��g��=�{��i�3�g�a/�a�Sh�8�,���K�����Q�q�9�o�0�1I12y0a�R�ʘژ��E�����Ù��173ϲбb�aqc�bIa�d�fYaec�e5c�g�ƚ���ur/��C{��z콸7mcl`6!66(��t�:�/��������ؿ�ۻOa�;�})�j��p�9qr�q�s�ptq�������u����8NN-Nggg''�K�K��u���k����0�I�P��uܳ<�<�<P���>^
�ü��i�M�+|������=�q@���jL��k�������O���Hx+�� �����tp]PT�Z�`��������m��B߄��M���	��Љ��x�$�4����=t�P��IQNQC�p�<�1F1�X���qjqq�����{N9�,A!�$�#�@����#�#O�tK2HjK�H�I�JqHK��*����v��)� M�Q��I���+{B��l��w��rP��yFy}y�|�����L�B�"����e�׊�J�JAJ�JS��ʮ����U�U�U��4�R�SŨ�P]SSRC���-�K���s�'���M?:�!���XcDS@�U��� ���YKH�C+SkB[\�W;_{��̱�c��p:j:�:/u���1�����Y����������f�ha��8�q��7�w�Bs��P>y�����=��Ƈ����L(LN��201E���f�f���E�ͫOR�4?�r򫅬��K6K�\�U�cV�V��b�h��6�6�lrlp���	�#v�v�v��}�+hl2V��8~9�x*�T���S��;gng?�f7�g�T�����nfnO�V�����@��3Z�=�`�؄��g�礗��-�)o�w������=�E�㾩�8�<N���+��w��D�E�o��a�� ��耑@��;�߂��2�A�N�(v�f�	-����I	�j�,�5�t��髧'���3"(#���<s��h�v��(P�{�k��"��Y��������}</s>����U�.��8v��R^4StPt�e�˩W(��\�tU��ݫ�����2���נ��_���|���)^)����]7!7�X��n��*�-p;����;�S���I#���w��޸�q��^gʱ��������=�x��P�aa*_jl*��ϣ���˞z��F���5�&�!C%#'�;36s3�5�m��6G9''�77>�"�7�*��@���P��qGQ�S�)��t�kqW�Q��g*�
��<�_�VS*;]��ܻ|�¾���D��*���j��_��쫉����XKĆcW^��}��j����7vo:ޞ|��Ψ��^��M�v�Q���;�w��UޗP�P֤�T�Q�c�'�Oe���-�-U�G[k� m��u��;;>t�v�vYw�t��������]��[�?;@53�2�8�;�dX|�hDi�fTw�����1���x��Ɨ�_�&N�O�L�M��ҟj�v��20�>=�:w^l����B�7�o_��߯-q-e-+,�^1_Z�_]���������ր��O��n�l$o�oV�D"��Z����>Q�&�/�K:�ϔ�&m��|J�b��<`"�-����)��thh��(��� `�M�}����PЂ� �y@
��5���C�(���T{�Ұ	����rB��N�p��ox��������o���^�*��Z*�_Lx�k���l ����.y�����ԭ���go���U<�ЇUՎ� mּ�}|CB�N�_��|�j��;�I�w�gdfe��>/-+���z[W����}GgWwOo�����S��+��kxV����T�����T�$�Y)�ٴO�ȹ��;'ts��cwy�b�W�:A����WI���.>)9��e���!J|�>���5m�|�Җ�K�ܷӟ���>I(f`���0�ﳌ��î$gW4�L�P5��9}�nN�ީ��j'|�c��V���������p�7_�]�^�^����e�2��b[vp��O`��2�Il�5�]�?i�����'�c� w��v��.�4��]�e��ؽk���� w����Gp������ ���?`�i!-�*�#u�VT�6�7a��tۋ�qj���پ�w�����i�7��R ܈v�F���;
ߓ�&���Mݴ�
�a(�w��
W�\cZw��(;��qr�Ry�X?P�Ogo x$��xQ��po�=� �E[��M����k�@Q���78ԐkF�s؋�T���ccSS��Wf��5K�(X�
��4>K��i�z����E�B���ٔ�a���ݸO�9��PD��}g��'��Uϯd^�Ј���>�T7���� EΏ�������3L���4���`R��	�w�
�R6Xd|u����ه�P�Iu��Z.��X<��ćl���Xw�H�#��F[�XB�Ʉ���^��U�C���fZ�>V��;.j�h|���K"0�+":?�#E�*a��6
�;I1jF���d1�
�/��K��ڷ$c/L�f�i��-���t)���C:^���[5�)�P�djK���:��������7�y�[x�q����5Ҕ+Ք�c�Yo��-B������Y�c�U f$c]��^QD=��;}0��A�/��F��w�,0]��m?��+t\tNr�9�0Y]|�OWN���8�/m��<����1�wW%�t�v�D��뮺|Ȓk��`o��� ���������o��O�W�j:�'��r��܎�����X#"�
|#�l��sAa�����HC\mMG���tl�����>m�Ec�r�}�Y��N'�*;n�|�z����fw���!��(���g�{��u`5Ӣ��X��O�dg�\�ܜto_W.�zϑ��b����3ň@�+���O�}M�	�Q}h��%k��Ր1dcT��fe�#4�}�&����(j�k]����{c-�gC0����b�~�_\�]���kT�ܚ|�y���+�Cˑ�^�Y)�_T֐3���W<<�1'�sx���jp�)_���;*n�؜��R*.wJ9����0���b���;뉊��J���	��p'6nmܙ�&|87��/��q1�%a^��]&F����᳤�2�3���%9����Yr�~��3�5���$_g�q��LJ7g}^�sR=)}h�hC1���6�Z D�b��b;(S���P�$X|U�C�����	,mƝr��r"�+q�5�,8}��;g�g��}k��\��*E�Aa��S�艮���,�ր�����v/�n�Dz>���*`�}|Ϸ1v�ύ��� �ڄ+��Tp�\�euP
Óa���Kv)��,5�;� Dsm���X���m���.l������	�i�ǻl�`a1)�Vť向3W��ۋ�I���\���mq5�=Ԭ��ܽq���o�Z�tn4׺�)�_�2�O��h:��� *q�%�Lʠ2��@���%.���=�U71!os���[�{D#W?��TP��՘q'>2?w�Т��0}j|��Zj*�.U�{��4�g/n�߶q2~�a�&���T��w���3e?��۟�ێ�Y ���<'�Ğ�����V���87Pϯ����:��yֱ@65v���e�^������͹>% '��v��7�A��.f�;�E-���P�/ݹ�v��=����KL:-�7��%ZܸL����m�mq��\����{L��rK�!"��K��}'�Uƈ�v5����<�lnn��G� �[�-�P�.GH�1��p���Z4}��9��"�"{���Vr)u��l�ޢ��jj���g+��=� �'�Q���G��K������D�Q̇�2�<4��9��s��LjSމ~�u��v1D��j�\�`9W���~��%�sz����N��_�?=���Fg����h��Jp��(�y�mx�=_��O���ی+��[����m��7O7\J����L(t���b&��j��8�R9��y�܀����������p�������Ƶ�k�� �uh�%k�pv���zZiW�7���|>��)�?��A9��K<OMPE/tQ<:Q��s�av�(������%�ÒZfYC?:��WV��Y.,��d����.9F��Ƚ�M>=&y�o�#�4KtW�!�ty��
}|<*R����̕�ە�V�Ӕf����̉�4L/��z\@G�x���]��U��_�P�=�c,1�el�|zA�k�姜3.8������Z���J�R��ϧ�B,9oSq�6AZ���'�f��kz�ȨJ~Y4��*�"�$�0�<>)��FQ�����u<ПQ��S/;Ʀ���k
�Y;l�:Wڢ$.)�dq-�(u��Pwv���5��ͷ��	��<k�B.Ô��ܪ��f���������g�5N��N્c|�=���e��_��o��S��.�BJ�t�iNum؀�'D.=�l�u8A��pq�[L���}+Y�>D�*����X���O��]�ԎX9Ӈ���v��.�!�E�ji�w��Kt�h�l��f'd��1�5����4�9[`0��d�![�I�<����|]ۜ��:/�n��,v����1�{�uz:w�_Ǿ��kV��:�V^�{��f#BquSs�y���6�Չ�'����5��1��w �m������+ͰJ4yח}�����p������cӮBV"��W�E-�z�|��ѫ��Iu�)�@$_�H��Գ�AG-͏�K�d��=yt���X0��X����f�b�|�hY^�Б���[Ny����% �b�U׎�BN�E�Qc�«�t�a����ګ���8���y���<5!�O��*��K���Κ�r�~2�o}��l;V��W��pL�/��h��?U����y:�r��(�������W*ON�z"*�[vQU��c�����/��>���>����7�F=X���_>���r�#�8�_c-k!36т�6Eh�K�:�:�}_�������<'GcN�j��~�s<sc�R���Uޥ��3n�<}�`i+�ZOu��u�QJ�}1����8G��a���Q����a�^�ɋ-萵aM&xtg��=+ɔ��x�{�ݨ�<]?���x�[��³ο+�{t!�.��:0��0���/���eo�brI�����m]�Df�ӕ/��|.=������k�/ß-9�����f����D7�s�,=�pO�J��\F�'���[��s����xT4Jek����V'�ݐ������Ig'D�%�ET���%��m���mJn��t���������"wv$��jF�f坫�	:���s��oG=�q=��[Ud�k���<Z�p�uo��b.�ʥ!-��8eљ��7�����cS�Q���;]u���sYk���qa6���"��}��oa>}<2�Y��}�׵Xl��D�Tq��<�!��4���0���������������UL�/VIT=��O�!GX��j�u��f�YM�P���a�}�XpZ$tr��� Q���oMxn��e��`o���fQ/�'ǒ����_ʺ�<G{GNL����sS��8�u(
vj��p�t0PAے���7�hmee��bu�R�@��S-���e��s9[2�*u8N�"�q�Ǐ��jm7���n�-�������6�<�ë�}����1�9�m�lu�|9���f_��;S�Uhӊ�6:�h�HQ){Y$�eQY�8�usZ��b�N�4|Vr�c�cꏄ�ULj[���N�uf�����4�r��6��X�����G�B�-�
\:��
i�. .���W[W��;n�B��n�P>�;ή�Rsh������lJ���ǆ(3V�D{v���S)���7�c�m?�����F��ޥ3��&�׋�Qf�~)�\��`uu�sP�̕��c�۾�/΂�C��l��2�>��P���9�5"p]����C�kmj�g�FN��֖_���& 1��Z�&�����(�ǖ?��2��wQC����9Jf����iy�ꀶ�z��?��'�v�x��UgN�8\@z�H|s�R�f~L`�����GSmW�Ǵ������M{F�(b���}B{n.�Q��^>�6M�R�28�$�����Z��۶=�3�W��+����u%G{i,�c����|���Dv�!na���hI���;���k�oCCy'�>��%F&�V%	�-(<O8��Ee~8�yh^��,G�h.W5�zr=��Q�`��o����n�R��c�=�/��dS�Y�DhT�L.O�7()���Tp~>���lp�j�~z��T��[���-�����R������U���5\F���E�,��4j���f���L�G���[��3t��>��������k��C�N���9UlT�!p�ýR�'H?l<�/���k�:���s��Ef$��N�q����`,� �f�Kj��_�tR����,��]�I��Ԕ�N���'��<M��.)8�~�-�÷~s�:�ԧ��!���c4���BI�}.�������,q�]������6i��U��A��i:|������U�%{^sxŲ��a�,آ�x���C�Qi�n�Xj���AXb$�S@v�%����AZ���ea����"�}s�33��yNiBZ�����	��=�e���#��r$��|i�����w�ա���������W{y��ʴǘQ�e�{�#�o�Rb��2�����Ͼ"���"�nm�Zu���kN
�ηA_��h.Y-'��� �x�fÙ}�5�ͮB���fx܇����U8����FH��j���)����	��ڷ7+Q��2�o7g�d�6��=X�sl�E0HK���c�T�+�#T����B�ofx��+R�~_�V5q���^�|�/��Q�n��o�6��e�:��{=�)-�Z���x��������n�f���M�2��7���cmb�Ϥ��s�P=���e�B��(ۊ�e���-�~�6�2�*1�y����$&[GO�v�؈q{�Z�7���e�Ñ�4�V6�_�S��g�@LЂ��g��{�(6�����x�-M]��(�"r�J�A�5gVHn{�3�0�+?�x�B�|����b�-TWt~;:��v�$��!և�n����o8�R���b����j�S�ʉ/��v<2a����	Qdi�!�$��f���3�>��C9$��k��Ι��[��G>��҉|U�?����|�P���63�ap8Zo��?²el�v�N���#�����=�:���IA*C+��$��c3ء�S7(,g�P\^�x2 �h?�Yӡ��	��Z��x��_��Ɲ���n�K+�Ŗ�c�D}��ךkH�%�+�^Pk\���J�死f�}�9���L�~��h�e�o�0��Tr�ߢJ���@����,�E�ߏ.��#��r������qӏ�]�J��m�8�����qF Ƅ��M��&��]`��x��ICm{�\<ݘ������\�
�#������8�άjx�P��dy�NF�v�a}u������
Z��NH":��h�zm�R\3���y�+E����=X6xEG���SڜZ0�����%���	�_2Gp긌����}�'��uQq�\ee��p�C<c�����S��o��֑��yqL)�#���i�'�c2����K��q���
��򡭥R���v7�+��͗�R� �֦�԰�Ȯ��6ܮt�&��s�A(fh�v5/
:���>��;���I��5��߈�W@}�>���������%ͼx{_��ϿDh���=�k�+���`���d�p���~}��?#{T4Jy����#Q�3i������N܈����B��4�vv�Զ�L��x�haB6�	@�t�'?���xd����_�I`���K7�44�q�Յ�'��]�!/��0WN�,�����yׄe���׊w��W݀V36;�2`^�#����v�fn����;׽���\>��_����e��zM�eܝ��;�yj���~ ��⸢��:�� /���{�2�`"�8iEf����G8�i�K����u�|�Eq�рh|���s�:</������������'�"���fȘ�J���ߦ�Ȯ���O?
�(Ǜ�z�e�z������ԣ~��y<��U"�-Q�4��+$T5.�Fh�}á�^k}c���̂�\\aűD��^竟�z�:~��o����WϢ�S��Ӝ������%��d:3|�	j�yػ�@�:�w�'�������+F�Z���|ɲN���������� �WB�G�Y=��ˍ��w�B�����ߍ�Z߼-��/>��� ����G��M�nd:��s�F�qɬ���Ӈh���WՔi����r��,l�*���MF���r��qVT��W:?��HX���c�p��[�Ċ�|xFy�<�h�4A�H�1B֥�W�*E�εܶ���k�x�9�ܓY*ģ;�mu���F /�C��7��M�)��˨��]��t ��e�P l���9��*�~������e�������f�m<�k�9�,O�S�R�����M��"��� �5���FC�9F�/L������X,o򭛾��_�^qI[&V�����CǛy�A���H\�Č��t�3ۛ�Y�:��`��z�d�%O%A�/�;��KZ"��	��#��'@��?��Dz3Ier�f�Y�&K0�k�O�S��)�*��������9�&Rܣ�ރ�t����S�>�lu�W� .�=�iK/6�4ov�=��A�Cʟ���F�\꾟�p�P2��՟�)5y�қ)��8��Y���+ڥ���ne�!|R���@�.���'5�٣� [���uus�aX��T�ll�B�%�_�/`�Q%� (^wtP?�$��[�֕w�wO��6%�ޠ_Z3_2�u���-�3e�	#r�3	k"s,���X_r�B���I���v��^�4P'�35��9����6טvEA��p����ֱ?���}��D4���*��16��6d49\��Y�����p���=mt��I@���xJ�I�C'MeK�{�s�V9H�I�a�$~B��^��K�̅���TV�J�Y_�ڱT�VM�N`�E�l�-]5X�� ��	 㵨y9�G�A��y�w#Z�%��A���(L��X��&4ś�M����N�������C�f�N�L��k� :�k~Eq|�M�u���ʒ	I<�
e5�A�뾙�g�����~f�����v��o�w�"�f�f��c�$W����3~�4�k����.��ש����b�����3]�Կ�*89E�B?L�㌍x��$a+❣�-q=n�?��!�2��{ehDFyd%1?�����o/�-܏f�rkl��F�$Uf�2�'e�~,d�&�.9�b<��u;�s���b9�c/+{����Jz��6I�O�u|:`N�Z��&KL�~v-���I��+MӋ��\���?S�_����0�!!ē9D]�?�`����7�:��8��E����w��t�!��ˋ%����p��`�N��퀥QBRQ�5��u>�st�}m�R��6y�@ Ae�)W"�+B1\�r��&Y��%��7Ԙ�-��͌ݳ�����ޘ'�d��m�ye�ު@��� o>�(�X��Dg�]_�G�(�1(�E��4i������y�=~/�C��� ���2&!{�m&��
�=���e�S�?Ӱ��5�bݸw~��[�A�#y�J��>\�U!�4�s�?(fO˝��o��:7�� 3K��J���;������Jd�h#h�B��p�Ў-����H+�H���}��z��sq����W�{^�F�s]>���,N����] � ���r9�b�����8�̔�@�*��`>t��8�ph��������&RB�4���Be�EE�ܱ��}�	�Ű�R:-R��O@X��R����R�2��cO��|Q�Ѻ��J�( /����7{�B\����97�^��rW}��?ef"�@�q�k�nLS�2⠚La� �̣ZR���!U�jY�CU����K�L}���A�D�wu��x�=�v�{�b��Ω�e#�v���͡�G4+��u>0�8F�"�sơ���ng�>����r8���3�\�MX�ś��>E&��0+��8��h��S��4�� \�@�F�����p߿n#�j+�y|qT���P�z>OO�B�,r��VKѱ���֥���	��wy9B]4�q��9�z����bv$'շ�pC�����
<����M�!)L��qsw�J��.�qWX%\�2pL��lj�'1hc��ŭҌ[���;i{)i�I?:N.�F32��7v�<�kF��P:y����ag��s~��g�ō1~�|o��a����Z�� r+q)A�J�w����<�����5�]�
��?�nǴ͚�
����^q��5�舆�4�Rg���x���m���R ���.�s/=7�@�%�ߔ�]O� �h�����z���`��UC֣g����;�~v⏧�Ҋ j���>E��z%L_3�*�7	�&hV�ބvob�吳g4��?�����̖�`�����[?H"��^H�lkp�_�l��t�7�J�!���}O�H�������-�����<N4�o2��m�#��=D��V��%��k�/'ߟ�h?����>�2"���
>�ւ�yb)����'ElX 쎥i�%z<�����浱�7�f��K?W�@L��n,�<�Cއu��rEw��H�QkkyC�OFvq��99t�����̓����4㭵Sq�z_�43qM�v�ʦ��p����7K�/\L������[��i�Q�m#�=\�����(XV����~B�e]��`삖���EW�kI͡s㒖��8��>��%1-5��k��.�7����nA��?�:y�s[{�� �g��LN�&��{q1�2�z�t?
??����/�o��:�ߩ���Z7�N�{yB&&�Qɴ����4�z�4*�/��5�k'g{��>kX$��e^3�Lޟ��<*��h��]C�fY�Qs��,Dv�u�l�TP��`��ʑ@��$ǃ�����R^7&u�n^p)Ki��7��]�3ο�o��J>��V�V��Ѿ���������3���Ao��QKD4�}��a�ѷ�,$G������׺i܈S�9M �z�d�8{Ӟ��`~��D)M��5�a��ϔP��{+���F��(��^�]=FD�Fě.'}X�� }1��nw3X��%�&k&��SE��+`~�X�T@���,H�*��~g�6ͦT<�,9��ya�T>�+�s.��M�}��kJ
Y%X�u��H�,#�	�,��7(.$$#�OU�c��v�xN����s�C�3�N⻙i�H�>l@o{�0Jt������n�YuI3XDD�l -/2يͤ����!yNiͭ����z!������ �p��x,��R�m��戋��2*Q�ڃn�������lL�J�a��n��oxKS�Ȇ�׆���N�G|�	0�T�$*H��4���D���Hۣ4�bf�>	�/��y�0�����9�����E*}���d�0�<���V�kx&�_p��� �R�D[��m'�`j�ϴ�nT`"�~�	��gnD�mGqXr�0_P�#�W?�Wս#��S�2<�����u?�K@F]�V�?x$�gG�x�k��X�g���H����۷tyֶ�$���γa���%���(=xm���n�[o��TdIK��l �MC�u���,�|�p�3�]���7�М$S28E9�d_%���ٓ���w�)�7#��Va�j�=��h��l)t+�O��b#�dNo�1�Hpz$��'\�E�����(�~ih�3	 ��Bu婕�4i��~ʶj���p��6���]��~X����G����!���0{��9�.eD�?�W0�M_7� �C��m#���`+���=�c��J�6Fa��jT|�
Sc���xa��;��{���c�L	=9��x�7b���`�^�sh�z�ь��g:Dj���$��4dF��4ٯ,.�aJ�k`�H�WG`�7ߡT�����Τ�=�ZtO���#>R�X���xh&0�ϦA�MW;���Ɗ|�~���0J/	��E�?������z�ZSu���\���}����3��\\N�I�/[�17c2C��	8f	�Y���;ǡȢ( ��R��1C��x���<N��룒ϫ�ʠ�x;�<<�L��_���k������|h���TgmO��jBL$p�%��	�~lIej�D؂��W��Vmk�R�M?E�"�	��K�W+�n+��;1�N9�WR6b����J,�_Y�
(���g�J���Ku�*p*� ��Ks>�p;^0Y-C�58|�����"ZX�د�����*�?��x�9��(T�+�<��=}6��ڧsLT����'�)-�ɠ%�I�y�2F,��s���=����$U��VϳX��>x9���+%p[dX�f蕼��BRFD6'c�p�������ްA2�ԩu���%���Viڏ��Z��R�;���k��]䳥��>B�	5p����,���E�w>=���ve��k"���n��	P
�f��'�T�<�/�G����\�4|Z��m�����٪6����6v|�h�C�R�m�=��[��V@��Nâ�E��,�	��9�k�c��Q\6(�^vӸ�|)#@�<+W�ag�X��3*'T�z2��#���,���5&<�<z�u���y'� ����}��iV���Y ]فP���*�zX�5�5�T/>��k��k�{B���F�/i���������'ts�����~<���g���������a�IIR���&�-Dy��qL
G��M$�v>Z�`����j��c�nu�&ur��ݒ_3	h ÝP$"2Tj����i�ݪb��Mn0*�\��B��5�(����2k��i����f��_jR
��c�V��&���$����(�}_]L�$++�/Hc)Y�ƗPV�'��KU�Iv9X�1챁&Ϲ�CƉ��z�f�ncv=�̺7��l�!�r2��I�M��{��'��y���g ���b���)�*Pu4ٟ���Ty-�RH7��D���\*�ʃ"ӷI�69�`RV����uaGg^g������t����pZ���A%6�:T�����/d����i���߈�$)��i���ݤ��}q���%Ͽ���3��f{�P�1�2`�@�V���j
�[����`�Iw~�"!����ߡ�NN2�7�;�f&"���~O|"���X�3�?��ڻ��f�h2҇�O)b>�r�%��
���W@RM�?<�΅�kB�K�����x��� }��ߨ�Kj^x�E]�q�$<�!� O��ʄ��%��i���q���w��p+�w
(E�e�ijw?��q�t���x��^:B����?�AY*W�],_��X���R2=��O�_!R���>�:#U(-ggxA��ʳC�2L1O�g�^1P�jQ|#���*T��m]ntݻKق�ݤ�޴��X������LX�	�K���nG�n��4 >�Cj�%ׄ?D�f�J�7�5���g��x��)���l	��qkG���p�b���-��@�k.tڦ��r�����t��lJI*(��f�g�$@{�,u����E�ƛ@|��;���e/�1���l=���=�8>T�z`�BfEf�K�����*�Xu6V=e|ghm���r�x���kH��Y�y�s�&��AC��2���g
漈b���ļ�G;��;��K	9���ov���Os�|�D�Xs&���VI������Ɵ�N����َ �x�-s���Z��AEk�[�(��l	鎄5�@�A3*��f�a�݉���uy�Q�/��>G�<�"��[?ni/N�T)����Z,3����i�H��*��v�"����{��x'W8	���P#K�R�w��Y���x&YH>��j�L�2�x3/����XZ1��TqT�̫f�5�E;��N�N��-Y�iP��H�u����&��ap���:����~N'4N�%0�I�ר���&�ܷ���]c�����[]����T���L�ѳ�<����*F�9��
��O�0�' o��4��D��U�)�	sv�Ab'�Wgy:(������ucn�<����gk�T���^�|,��������A'��^l����$5v��[[6��C�R��L�G܋T��55�-!�0?�wՠo�=cy��A%�<��ܡN�.�Y6U�\�׽8Z%���eM��Y��vтX�	_#��2�_up�zȇ� �ۋ���F�Fę��T{������`]�!@�SrW��i��n_s��g4���W�<���4��~Vy�F�R����"*Y(鹎��N\"Û∑!/�L�$i�7�c�'�ov��\�$A�Ȍ��'UO��OO7�,S]�*;�- 悰�n]E���PW�d{]锋I;�c.�	m3����H�m�
�;k�'Zf�B�;I�����~� �p�����f��6��ܝ��Hk"��!���@�
�����c[�?�v�s��Mr�L�z���;��3J��R�ʱ�.��*�z��]g�l`Y���"Vu,�2d�nl�k��-�&����?w����k�eK�4�������e��D(��W��r���<�楈�W���&��v�iqMD��v`�r�KJK�5�Q<;�7,MO�L%���&���޼��Z^���~�+J֕�*@�f��ѻ��nZ@o�nr7x�u�Z���Q���@C+ҤRlG�Q���R��]'��m�-(��ׁY��� �|N	S�U�1&5�J:{��i���eU��֕�S#~��|�^z�᣷Hjhz�;��.0c��Q���+#7��DE�keN�ꯍw�9�@�*VF����U�Ga+�ҽ���d�7�ȯ�����r�w�]���s|�_uNnW��ΐ]�Vc~����X�2�3�"U��n�� �\��A�a2��"g^U�J�ȘʒO,]*os*"���\�#��!����C�]d�e\47����Zp��;3p���<%�%�Q��Ir��k;�+���P6��||�:�h.q�ޡw��W���L[ĎW�wN��������ֵ63}r֞�A<�.�/��4��e�q������{m	:�,���l\�3��NU���kP�&~h�RM۸x��5~G����E�o
��qm���v���Y4]�%�k�>{0�-�"%���h^�	�l���q�\h���
�4sso�����>WgԲ��Dm��=��s\Ӣ�c��,׏�1�׆����,�%Y����S�.��v�_�>��i�>BG���E��m�Ϋ��	`���xm����K���*��U��T���1r�L��&bL����5�9+%g��V�*��~���l	Q����0s�p)f��֘x�Y̳"n1x�mh�u�zْ��ƇKB�2f����ԍ�w\�HRX��ڮ�7$�6DNAvJ�Jk�$'�#A<�hŜ�x�B�)>�ޞ0�|�UWK�hw`��q����'�G[>�WѨ��Q�uF�N#���}�U�r�t��D�J��"����p��0�"�"�x1����{��h � 0���tv������m����֒ijH��>�*!�j��U��ϼV�iR�9A�i�{ErUx-Ǥ�$�(��?�����otl>{OtՆ�{�����|q�������>m��d>�`�C�Aa��PS��G�3[����(w�
ļ�,ϸ�^W�Ԁ*�s+�gj^�a�g��ٴ��zK���u���u�u�du�����^�U �� �Fk�=�dRRw�#�Pu���V��W,�.}M
nq���2���N�����r�r�i��{Y�����>�����,n�v�⵲g)��>`���=L�����������H�����T�ǅ/�@N˺=Ӱ7��ޱy汋�����T����B`�c6��AŅǲ%Z����hH��0�6�,�8��h�X�k��gE��~�f�x?��!�zc��A�Ll�q�[2(Ж������"��b�9�N��<� ���XT��@D�>���TT627����@4��궦#��+�n���0�3����B���|���7]��Y��.[���x����#2��A�_[�+��<>��y������r��C���0�.��u�I;�TcZtd���<��/i7�~,�V�M]���[����]4IPO�.��o2��WQֳ��{Y$����(������TAC������rt��G}0��:П6g�V
!�=1:��Š�Q�1�����\Y���p�F�S�-���jfUݣx\_0�3��<���k�Hٳ2���5� 1M0M`-ѕ4#G[����uu�_4�/u�D}�u5�	Q*�_����>��8i�PL���_G�զ`����ƃZ{l&=�w+@zQ�+�^?���+�x�7*3]r��"�5eR+s)G?������Vd`z
X�Q�(�%�Ua��b���~8�e8��xI9?�\o�#McY0m��*{�� -��L8^Gv�����d�h�����Y<���F�����fT(;�jfe��%\9��VLl���3���v�0L �1�%T����:9=�N�\��w�~�N�s�%�Q ҥ=�諽z\���t��l�L�����]b�y�D�9����������ZT�y���܈Ag�Y���'��+���ۊ��u�ǈ?9�z ���vvy������Z�6��z�hKbE%�WSQ*Mu�f���}���;[Bwئ����ݓ�'����o<C��xʋ�6�R��#�`v��
Ȃ��4"�+G�S%��L������a���L,�ѳ' �h���!�9�~���D[t�q񷨲C����N4&���>�]�������`���6�A��E����`|[����W��9,�/)��D���p6�YJw+RA>L�*�!y�5������Tb������,�)�/=m��`8��� PV>l�p�v+}�����(�u��X�C�Q-���%�BO�O5pq\	���{�ز�����9`0Vr��������_�q��>��n"g˗�J���-q�K�Nm"��қ�o����7�?����� �ڡe?3��Ԧ3�;v��J��dhδ��c��N�R�� m�kVL��+_��%
��y��� � wל�Z7����H�4�����'�����K��j%=:ts�t��w�^�v�P�B�ޜ�(K��w��� �Sq�;"����p�(;>
:���zw���Cf\�Kz�HqǬ!	?�Kq��	�K}�bc��p�t�Uʳ���"�DQ�l���p�0`I9�J}��G'Ya����X�a����k���}y�}2���K�v��FwO�_�As[���?���V�6'�C\�t��xg�,7����c2	:8|�R��8��Ĳ�a�#G���[���p��K�rr���	ډ�RI�kZ�D�v��^�
sdP�r��V����;�@�H]�zj9�*i��o]Η �7�i5C��Z8>���@B���J�b�4i�{�K�5�鉱rYc~���R"����79�:��t-�ݾ�oyz�r2�oe���m!��|)l����e/,����}λ���#C-�v ��T���V�]HSx4�c.�r�x��1����6Ŏ"jm(dw�D�Hz-R+��FIKK[���1��h?f��r�Ş�1�}y��R`>�߹ƍ"�ȗ��_k!d���NX{K�B��,����ռBw�~�y��/��>�=��m�"�_br�]@]�$�����T���-�|�o�i�ޥ�YhiӸش��$O)�骽W7f'fd�\�y�du�Q�s-�(���(��#!*2��͹�qi��|��^��ٝ(qc �a��Gm��������ɍ�Ҷ�#A���$���n����eC�9��������&��Π��<+D�t4��"��c�����*�4��G��t��������e# �F$�v�U<�q�$��x_�d�~=t���CZ�yT��X��9�hyRA`�911�^_�u���v��=T�S��q�ܐ���!��-��Y{t�U�/������l�piZJ
m�Q�����+����s���S�1�����
ݏn¸~�{3�K-k��	P��-�����2]���fO ytÍaǜ���X���Lu�������f����O�:M����x9`3���;ʈ��J�S��	1|'Q.�8����f��8.g�?�b�����u8R�_�T��2�x��"�?E>ɻh֘�o|Lk�06�1޹�69��`L쁩����95����	b�p�رH�K+y�pAy"h��y=/�mi�"���]V��52�E��ʾ�;�����S�]��J����;��ͻ�Qa�����s�/�o�5�)�u�WQ��ڒX��YFX��Q�^m�Gs
�M�3��]lA�x���͞۞�T^�m��u��㝆�+�m"���¢+��Ψ�/��hQ(� EJоa�ڇ��g�0���1h]�Zfl8hx�[����Pj�� �)�J��������ޜd;�%	"�Ӽ!�j,�\��nϛ�[�:Ĝ�n�_��Mx܍��&�X%�/㦖�R$m�j� �U+4]�����W�?Oj�T�%���8�̋��`~�2�v|I�*:���r�5,���4~/���n����[�l�u�=�)�ʆF����@�}����̪�vߣ�>=y��F�`^�n\Ix%��<a�F�D�Y2�S1�CW����B���Ǫ��Z�+7kW8�Z%`��1�Ƙ�)k�(�����PObJ%�2G̨�;�Cŕ�0���Q4TDŧҗ���9{S������nc�f�R;¥���=4�����D�p�.�$�>�*#��� �]�:��9�.���y�(54�hP^�Hö�_��Q:\�O�3�y,_�R��]3�d��g�	�������20�Sk��^�"�>^8����7�SzE����N��=��4�X٤~}6]E���".7�4�[\]Vl�Ԣ���]��7��*�g���c�$�ךs5@SFǚk_e�����ܶy�x�B;��u5�����S�Ӎ&���+�{vU@��X=�wQl�T���n��o�~�9�+ O�6"%����??����y��մ�����_!�y�,�~~Զ��;�"\�	-$zn<�G�1X�M]���M���	@��3P}������@}9���V6���;k��M9fj���,������|�_0��ZZ���"�~@����d%$Xͯ-���b���T~���o�GJ�{WZ�h
�?�� \O��*OdL��� B t�WR.4"w&�^;�!j]���r*3�t�]�TKr�8>�=o�@�W<�Zd�����t0���k���=�ajOӕwͿ��e��|�3hq��o%�V6��tt�E^��~�y>����DRz%��x'�xy���@�?�k����I��6�=�p�N������I���R#R7CF��$�p/dz���ԙхx �ޛ�x,�{��H�'e�A��0K�!�w'�Y������$nh�ze{��sߦ(���l{%���АQ��o^�+����4V�L��|$�)��=o#2ʋ�����i4+�:,n^��V%;�O���Y?�|���ms���h1����֌�%S�m�[��܄!�9觪�-%O�]K(��ǒ�p�=E�̚����S7F�A�8��咬��lr��vЀ�ί�'k�b�J}F^%�,���D��Oњ:L`���%�~�nxZv;�P��?7���f}���:�M�Dd�<z�Z��+����K�q+ٕ���,H��;{����.�C�EMC�1q�	�s�L,���=�Ņ�9�fm���R�$;��:ş��b-�\^�o4���\4b���M�w}���`K��u��PVr�n˔$�S�u���y����'�Ie���Mj�\�����F�!!�(�W]..��@�$y'^�pu��E�#rg1K����bu��9$��ٕW��P���/_�v���ԏ���$<�A�bY[��Ɓ?yYX�.5�IY��:�bڥګ�XQ�ǳ=BK��ND\Q��L��/��SS8	 VZ�<�b�N$~x�]D�6X�Ф	��fH̍���0p�ZY�;n����?��9;���6�Ascg�kB����?\/i�΃�o�HX����-�Xp�C�Po_�C��>B楇�ī�$b~��-J��u�'@�޼�D#��?���k9>�`�%�L�ʔz����^�7$��"Ц��T�<Jx�~8b!��0�]�B^5�F9z��:���������*��;�К0��S)���Ұ�ePmg��!�3�f˧\��s�xW/{�o�b|�W��nKW�|z5������J~�P���s8��Q��C2-gW���+j˜wn�yX����ڈ���S�n������~5zY���+�_d�Z�u{��cv.��0��wM�-d���n�[٥�.�HI�hW�[�kA���@h���V#Ƈ7���t����Ր�C���MGӠ5�� ����.],$��#���*��A�޷9obj>�IP��S{B�R�ug*����u�X����%8��B%�-����a9ʱ�R鴩��<:-��N*ƹ�/�4�����%o�;˗�45���[��S��kZ��K��+��z={�ƻ�2+~Zhc�+6���GY������������%Mƨ�Y �j�mBX�}�O�=5U������/O�o-���ْ&���0����r'�7�\�Z�Okx^��;�r���zAܰg�|��
�,��&���8p?}�D��]�v�J�q�h�c&f[+���*K��LFq�r����iwzߍ���Z���R{П'�[�dh�n`K�2��_���a!L����jI�L���ွ�@�v<*����3>�Dڜ|g����'�߹S���J���-R�{�$�5��Jʼ�n�r7V$��$�{�m���}��ku���QVQI��\ݬ>��t�
Y�.�+o:{���@����Aȥ����7�j���~�����QA�F1t�ot95��������!�Y���ޏ�2Iq�;5��J�eX^G�N���-��߻/��� ��L%2���y��T�ſT|y,��Q?^/����>4������-��h4���\G��*}�xk�l�䈽D�K���Ȏ}�N�ԕ�4Ja��<�V�v�8HB��3��J�Xz��#}�/�at+OU�Ri	������Mb�#�(%8��pvm�[�
W�򭂅tAn�a"���Z�kǬH���؞&������Ta �K��g�Nqvպ���[9�*j�
���U}/e�4�1��oɩ, ��L��8Ũyy�mR�x����<�g�6���6' t2-J۰��C'��v�[�����/x���)J��b�w{���h�y󶛶O�jٶ#H�*��ě�������F�X�����t��<N'�նo����T��&IP�oȐ�:ȹ�t�>۷����q��/ʦ�h5��I�!x=�3�q
����.�b7���F���Z}j�k��C�g��%�seD�Ǟ��&��L��g�u��\. �N>�U�|s1`�>��JS9[[�hi���@�v��3��Rj�ɥ�&�l�������$m�K^s��y�TФ��������~�)��JrV~���U])�x�,`��S���-�I�o�vE�Ԇ�G^��QHif&�1!�>�����6e��_*,k IW�T��վ�Ǹ��i��ʢ:��A#
^$:��[ﶈ_� ����h-@�����q�=�X������+�n�VV��%��6[6�b6Y�?��l��C*��Ê����u�h�4*
(���Q{g�J��J����J���>�z7 ��Km��Bw8�r9�	Bʁ��/��a4�bȩ�zG5q�p����OQKʔX�O^�e�֕�P�G�+2�W�<����+/95���of98�����=g˄_["��1БF���F����f~��^����%���F/9.��t��		�E�BD��sQ��)B��o�[n��F���v`����~����[� 2 ^>�V�
���*�Y�=pl6x�}��P����ܚ�go�q.���-^�ה<�F�=4ãz���X�2�\����Bb>gվ�9eX�x����������1�Ug�w�b������G� 6��:��,�m>8����\�c\?ڲ@"�l�Q}�e�	˨D�'t�va8ƻK���y���8�]A��^�/�x��7�4�R���^_�_ ��j� �FG�Q!/���i��V/����)j.o���b����n�Jl�2��W1Q��.��/7P�_�^>��?\v���]����]�u�ә�N[;�k�^�{��{�7>� �J�|rš���O״��Ð��ߦ�6�<�#�I5_�U�]	�6�.]�š���ֹt�E�� Wb^2�t�7w�+""�J��l�^�(���$˽������	!�_�P�k����F��i%�H���o'��S.�+�ߩԓg�I\y�1�����\^�:Ϣ��[�$�5�AY�;��d���Џ2炧k+V7D�N�%�Ln
06�lrm\2O��=pc��w�kÖ�#���[[\]v�-���}��<c��;3�7m�Q��$�AU�P����͈G����d]~f�ܘb~J~v�D��#�ǫ߮�cq���=J#�X!!�4���D$�;�z�E-ѡʝ��ԁ���l��U����J��F����j�{8��$qSR�E+/�<&o�%�ˤ��Q�#��?����g>���wܚ��-�F?NW1gf*����~����@��W�F-YԬB8���.F������i.l4	<�b�Zh��*+���j�?̝u[\��i	�S���s�@�C:QB����[��.iz(x��~�s>��Ǿ�Z��Z{ߛ�k��l�"9�3O�}�g��N�6��uU�v��"|w�@�����߃�ŲK��Qc�F��U�h�64�������{,��㶵z-�4r>Q��{h�ӟ�V�f�E�fn?�^��bMD��s�ɯ"��L{Nk����be�i�>,�*	[$�Q���e�Âj$Z�[����.�ߖ�r��$�^���V���'Y@l9�Mg�����;u<[<EM�~T�L�U�������{-g�ib��=>��Qb\�SX}���L<�t�!�[�����]-7�l�	f���nY��C�<؇��Ob���؀�" ��)�iBq&v^�b�'*�G?�2"��#S����g�s�z8p�|1�%-{��<����2Zi8�DK2�����(��	*]����(���	1�C���v ��?����F�H�Ԓ|ժ%&х��,"ӧ���]f�;�e�옋*n�#�'_�$A�d�M�c�B��'���"��'^�:"�:�V;�x"�����B��JZ���۹>�FaU�8�꒛/��	̀r��L�C���6�z6n9��'HZ�2H���-	*��J�9�1|,ԉz~�N��0�زݿ�+o��Rr${�*���z�ߝk���#�ħ�.P�t����gV��9�2���ZĻ۹�~�C�t�T��n�LiK$i�������YV�*Uqt�M�]f�U���k����߿b�1%�A��g'�~��Qy�f�}oC�P��(WC�v�C#ZQ'^�e!�x�u(L���lJI=�����ݶ9�ETp	N�!��w�Z�+�#F�Q�}��I]�uh��O��R���0��\��c+�*c+�֜��'yh��H��pejk�����E�9:�.��89�:d�*2Љ޴=���t�*%�vQ(�M%}$d��欻J�	jR�������X}�#�\P������d��>a�]�8n^���n0��,-�P?�i�8[h���cE�g>Y�u��ܯ�J��w?v�ڛ\�r�i� ��P��Z���u���yiK�J�(��BC��s|���Nj
�R/!S(�5����6Q[�bB~�l�kP��7H��|إ�i���"�vc�i'F��ȶ8�ԫ�~H�L���j\�*
����T%s�~E���d�(WmM�&7�����,���m�(*ݻ�y"����y�d��yÁ�l�AG��4A1U7�ϴz��;JnO຿�ɍv��5��h��R)�f���f���Y���Y�<��K�s�aA,\n���c�9%0f���癱g&�;/���ι�=~��>�=���jn����/��6����9��/w�|�I��O���5]#���
Q���=Fq���9:E�@8\�c��{�hh�B���E��!�K1�t�@�:k�=*.���iuu$9;OdD�s���ܭ�Ѵ�Q��������-��"���]l���"�Tz�G�p���=_p�ޫ/헟$`,�(z�6r[��s��ޫ��5��)R�-�#Q�	g�L��4�N�K��g�VߵR5��_��崘����Om��H��Z��Z�� �)��H�U���G�t��ش��w��!;f�`�V:�m� ���pd�1�T��J N{�����'6��x%��'9\��4�q��tLg��ҷ�_.�2i���s2�w��V� ���ۨ>J}"�����,���+<D|]H�.0�ĦWͮ�٫粬K�Do��4��ۗ���ݣn�̘�j
H��)_�%���_�`Pd�9�aD�,��z�Å(�����x8Bs�V�9�Ѷ�� &���Ha�{��.T|O���
=�b��}S����&��Õũ8����_@�,R01�%/.�N'O����oi���/_���S�MUp׿Xl^6@R�a�p��L����i����&Z����D��.���$R�����3�&T*�p�.X�N���vj����6��8)#A�n�r�\5�71�;Q[c��=ⲋ}p>������}�%�������xɒӃw��1}t������԰��th"���I"-3ak{M��B����@Q���Rs-2�d�e����l�B�װ���B{�V���/j@h��ft��X����?~�Ex�W�՞0�f��jfT�p'[�`��=�q>��!�o�,��FLM�
�]��K�ז��rji���&��|z4I9�����!=j0O'S��{\]�]H ��+�����3f�&�v��� :e8Վ@�O0[YnY[b�nFDh]����!Բ��p���#�����CMzB�!�c[���gЌo�Ů�h�tf�>���q3 N.m���֡A��I�'���Sa�_�)�������7���K��$w�R����$f5mr�?q���x�wD�S���O���X2���AX|;)��ݦ���Tw��6'�I��ҶF=Y�:��=���z ���wq���zL�6����7�B��p��Ƕ;���
���Ț
H`A�X��Ϧ'��,�V���(�--����l.����>jK�`���҆x�J(S<
�L��f��-�ؿপ�U�g�bmԙi�|�L��';�{�YU�Q��pr���)�f�Km��	�J��p���b���Sοk����\�|O��FF1h8��u�7�?�7�q)�}�[��ƺy�AB�ܚ�F��]��͇L2�+ cv;2>%�v��o]E���M"T�훶�G�di� c��Hkv���y�(V5����x��T��1w�n{�j)ob� ��&��GMS�F?C���؂����b�/*�Y�8��>�K���ΗB��P�Y�Ꮵ�����<��-��� �>���,Hܣi�7U�O]�?�k�����H{��$��$�Z9b�	8��-Btۃ������0g��e� ��:)���σw��!��W�G.��pcj_�隠'�x��Fm���ސ�@�ߥ��A����V�5C%��Ɵ�OR�k" ��r.?/��5y.�.�Τ[�9Z9Ҋȸ��D2;�eu���C�$��X�Dp�B&O����+�a��e@mֺ��� ��k0y7J����u���Ĩ����hzY]�'��,N|N�Hm���%̜$�-��#l0��x��z�/��kKM.�����y���-sEq:7Ѫ���BM�� Ĭ�!>1pܹ��R�%@����4ֶs�r��ޚ�@�J,#�a2Xpͫ=\C�U�B�Ά�3����b��|~b$��	�W���I�Һ"Σ�%N���>?�z��T]ĦR�6ٟЏ��'M:1#�$��L�q�W�3bH���"��`�S{�>�C(��X�V�������{m�1 �n��.߄��-��!�������m��E��yw�r(�.���/-�ؖ��ӑ����1���>����1���h�	b}��%�/��%� �
d��z�Wiz~�/�Ǵi�+%�8�k��!��1��	4?X<Cb��yӈ<�������K��/��Nts)�^�����T�/�2-6\n�[� 
��H����?F��Y��J.Z���-?7!�o��gj:���SK-ۢ�:�h���?w�^Yߔ}�}S��S8}s*;u���^����(o�Y��#�c&�T1}K�RG��W��m�o9^�A��fjJ��KZ�~����g�5HB���������v5� �.`:�eѐ� ��^�R��eM�X�l�d΋p�_�~$m����o
�������c�A�+��BA�-�/`0{�;���yCu�Uz <������7pzf�z��.��oe�բQ�eh�z�,C!��������>���0z����n��(�����rU｛iK�����x���c)&��F���V�qOͿ˺z
��uq�z�J$��~����	��_�^.���i��l�w<�cg���o���%���A�����J��]��/)b�:��������͍�i]=\��a��$��L,4�܉$)����}4�Ѷv������w�uw7/��
��G��'x�/��2��*f�he4�Wl?� ׵$�j����k%)�q�O�m1Qɵn=j�f�6�'�/�q�&���7�Tͫs�Թ�A����J�i#����{�x��oK4�I�>EZ�n�5yS�"�P	C�?WVyC�5ذ*��Gz����y����|tC��#���,��uje]>_M�j��N9��Z�;��1����! ������2`��ǥH<T{��ᣙ��}�<í$-G�l���u�7����1Og5ӗ��u�ɻz��=�����o��d1�櫘U��I���������~�V�����h�a�y���s�s�AԪ�y��Ng�16�9_��l.�������S�Bo���ar�"�Al�A%Rj��a��^uK��<\�-��_� Ƴ��h�+ kY����g���o	�m���Q[y�i,�����Ӫ���r̖�eY��ӂ:>x���� 5n�Ʋ���%Q~�9�PL�u6�b���S�:(�T�#��=�f�t�J�	LL?��0��SC�"������Jq?*�Ҕ��<�]�>yB�B��l��`e6�?c;ԅ��_]1�I^x���ݠ�m�Ӱ�$��#狲������v�'��5g(��4�x�%���e����s���+@�8p�p�t+��|��N�$���L��9P�3��\~�G]k����{�dƈ-s˔a��������ɪr2I�񪢝�ӝ��7���p��s���Һ������}��>�8zi�����w�
\r53Q*ÖD<>b L��.����D�{\F�TJ�__1�=�N�w{-�Qɼѱx�T��%P�e5ױ���^�mH���FLS����3�}��#�pd^o��]�F��1˱�As�-�%�'s�7
�،@d>tߊ��%�<h�7�х�=�3�a3����W7%_�!C����$V"����%�%��w���M��*;�'m��u���O���s���%����u��S�m���a}� ��`P<��M>���}
�@u��`k��D�8�T�_|��嬘����r��uᤏk\.X��pL�Ŏ���ET!޾V�_E�i�ݪ��n&�����.ѽ!�J@].T���-c)9�X�P�? D}/�O�=[�yo�i�
7���˻�N�M'��),av4�ft����'��V��m�}��T� �F.��n������E��������F����RG	���Q4�����K�3_v<�<\=�h���M�ٹ�`R5d[�8�S�UW��~�� �#o�}�:�Ξ��]x-�7[�<��s��=�������	)lQx	9�H���ܜqU�`z	�.r>b��P�y9t�q��W]]���(��+��4�P���tU�D��Z�,II@?��"�1\�q�ϧ5
���pL}�$c�_�ѿw$p�=�i�v6=^M���(J9}��p��K�w�#��̾���g���I������ݟU�M�*�},0�!�r��������G�
�Q���?, ��*��µ�D/'�+Ad@K��͈�V����YPh����0FuL�/���V����d&K-HVC��J|{��Bu�X�
`�Nl6��yX�:���蘸guw�M�HF���T�Y7=W%���T�6~()}��:��ӫ��7ԝi$0��$���;~�p~�̶�)^�O�f�6�'}�)($�p:G4�`:�C�ٰ����G��۝~8�ݭ��T�&"���c��
�-f)�-[+MD.����L�L)��ra���+Б)���ҁV�.El�ͥӕg�M+�-�Dě�u���*���k�����jd�W�s�v�,l>œ��e�͑$�m*^y� ~)<3N��Y��L0��"�����(�ԓ�O��f���^�f���3�k1*��� �̊2߱�����9)e�
f��0�`"�oִ7����n�E�D8��*�����o��i��<����j��AIh]o|�Ny͋�8�a!�����SLS�\?g!l���ק�ڱ�&FI�7�*L B7���'����ɖ�1!�X�|��|j.f	[KW����I���(C��6_���A`��݄�#%]0�)�N}�fD3�g[�]������e�C�F����u<�ny��6];^ޘN����=�F0��_-���`B�Y�χ����\�GQn��K��^nX�hkÓ���:���"�޼=fj�x���-���4�7Bje@�x���Ε�iobV��p�\N���/�'�j�&��*O*��L6��F����ؑ��_ߴ�5�u���pؤF^)����M����Ĺ��=t�'Ap{�R_�˘�S��(�I"di���������©�bh`�)�s�t�ef~���8��'�M��\�}\w�L�/
ڄ���M��`��T��t@}��I�!mV����X���ÈZ]�P��n�@N�9 �=�d(�]��:	+�G�H��ӈ��O/wZTHңF�	��Zlwʤ�؇f�?�����/F��n/QM�������ڹ�Ϳt>i)J�,��ϙ�X�)'�,����I^���|����0�^�x�{�l�!���hڦ��@�H�Q�Xf\`�����؀joc<����3hIhAKZ����NMMTK����|'$�-(�Vr��7]��?�C��y�S��"6]�ެ��Bf�Q&���W�b��0+��J`�C�/��gQ�D(��a�O����})���G'K
f,E5���ƞ��UT��*�~մ׼���W��o��<i��\���M��R5�C�<#�ϳFo��X��юN.��<��v��[=�
M&2\)Mv��~{5�g��q?l�����K.V}&d�S22.�q3Z�UՔ���� 1Z���;+��?��E�J���g�M%a��'	��K���>�����[�W�s�"o=�P'%��F�i�Q�oQ!,��|D�#�`��%f�6tb�#��Ũ���~�~-�i�P��s?�e�=�o]��j���1dR�/��S���!���t)Ȏ�m��]�8��4�C�_��z7{�}k>��B�G�*3������`2|~� ���.{��t���ⰴl`��Z�~Q�m�������ч洸k�&�D�E��wڇd@u�J*�@/a�-�|^�X9����~zx���.a����)�[��&�N�o u�s�%�i�ؾ���Z�x�pwK�i͚x61�i��M�&q��aaZ���ǧ�����!� ���r��xrbY�{��n��R����l��b/i�,�Tq�����:T�qM�d�e�{}=ҷ��2TC[���f׫ի��ϝ��~�hݟ��:�ڠ�H�2	�Q�H4���j�>�i�S=Yժ���������ņ�S��p�e�rn��n�rQxO�TK*�D��Q��Qb
@��`��_�J��J����6T�;\�W��d�<M���}pi����[��6�ȇj�h�ZW�|��2�b6|B_n��{�wl���@PrbO6`��G��T����߾yp��U�v�|=�U+W����b&�iϿK�L�{�w]������8Q|9�?�7{�){*B˒�0IH�f�[���ܭ�"�\����%Տ�"�w��ݻv���:64�I�KVK�M��b�a�;= �Aп��n7F��f�U��\I!}C�zT���-gT��f���(CM.�vo��_��|I��m�M���N�L���Q�ǉ��ڵC�~#���':�Nb�o6�%8T��*/^�⣸|7G�K��Wp��O-�[z�m�O~5�O�5T�P�Eٛ	'�-�P�H��!�_� V[�N��d=Hf�T�z�'��E��YUAr5��/����_�R5�?�Q�l�c@:�ڳ�~���Y����T�VL(
F�=�򞭩��b���ř����G�����g|D��iVf��̫���iJb�;"O��^;��e2����-ٸ灗]բ��y͖��!�j�''tƃ89J
4��12�1�ak���wp9��xZ�o�:'쩖�*��膺�0,&!;���i��Y���'�ݦ��ae��C���Zj�s�7��~*s8�����'Ƨ7!�j�@K�U�( Se��"�|��2u����4�%�?�W�t�(� B+zb�=�7G��6�,`	Dqb"����V��Hľ�;��%6z����fl�0}y[�l+�v�
��/��5�&�Qͧy���9�;m.$Fݎ�&$O,l2
�s+>4ٖQ
��P�;��&�_.1��T�|�6~�%�St���T#ܹ�iމBz�V�E���w��ܦ����y-`�3:�����/٪>��	��M���I<K��ji����h\�S��C#�F�?���ٖ*�}�@Kk�FO����YP7~<P��8����D�j�0S�3�[�
��^�C΃� \��^�D�-���T��|�j��	��'^ʷ~	{**��u$�
���/�N\e��"|>��5�7OSv]&-m�'�NF����C"D�����`�����hys[�����q�tjdC�y�I'��~uCD��,�!|n��n�_�u�(��/��C.��z]�_,�j[��P]A���7O�礰.q�i�d�������(y�D{L�F2�V��/��:D�;��%�=��_��r{�ߔ��|����Xc+�����H^>��������pFq_2�$A�Ї�-���|���(�a�i�>98������K����w!*	w�MJ�s4�ד$�S��#R�Q-�tz�2[����`�����F��m�<�C���Y�>�R�vO	�q�H�-�LT~o^�*���?,��,&򿺚^�?���|8�Z�Dq{�����_jS���i皛��&��)�`��`>u�r����9i��_O���I��K�&c�p(�h3�,=s�ѹ���i�t���!'l�@֎'���_ҫyn�h���j�"�7_�~2�Ȏk�+�B�����s]*6��?ɕ�/λ�����i�s��N��W@�wE�*8L����+ #����0rX��b1@�+��v����c0���Q��ʂFz&1�����/ޓ�Y��T���+��*�|hE{#��I���Y�zf�����P������ �]�@��̽aۻ���sŔڵ��'�v7^ln>��}�2n��Ê,���Q�'Q������/���|^!�
� ���}��>,�B�;j���F~g��X�x���&�˩�vB����v_M�����T�
h�,����֣�T��e�J^&�ߢ5ն��k�zA��A�����p��Ɵ�k��`����}��)A�t.�,L䉥KO.��1��{�}B���@kh�����G�M�p
]��+�jqz��W��(�֋X��:<GM?�ʊ�����a��)~�s������(�����`�ʵ�/5��#`�g3�~�P ������B��g�*��dycڿ?%�Z��j�����u׹�� mq��JW5�<{�j\�`�*��;M9L�d��:I����7�����Ú��������b=���Y�O��,i~�d��b�~�|{Z�d���!r�����02���j'IdI����KC	q�G>W�鄹k�o�>�Kr�',���%4��x���*Ir����{��I�b�L5i\l+>c��w�q�V�C}<&�4�rp)��U;� �z�|����n��Z��mVt#C�8���ھ0�`y�_xI�U�q��������jx��c��q�ɠJʳ����V�����VG5i�Xr��r���dB!���~���9��b���������T�sgܘY��]6�l�����N=z0�}���Sq��z��A� �v��*��7�]��� e�S��;-�J�cKʶ�R�l��e5��7$�����r�hT�S��f1L^l�o���y�~5�\*�N-�ynL�^���q���È{y�H�W�ްv�	����犆Ņ�i�`�s�\ލ�a�\���?~�I�.2:y��$b���з�Z���0��h᤮�}�/�I�_����$jJt���B���0g��ҕ懥����i�;g݇����Z4�������:N̛9wB�Z����$��ۺnVme�D#�K��E�G���%�&�E�1�h	^��h�D;s� 7��s'���aj�Et���&�֬Gſ�S�f�w���O��iǛOz�cä@��}�q���p��ȷ�T{�y�w��V�g��}���1���h�� �rzI&BQޫr�!�� �Z����a�O�oK*�^�����0�F*���߉�2V��k�ʌBG���+o�>g:'K��+�v�or�Bg=���=j��-?�iLw��$�
:�`�q��e�8���m��k'yS��e�+�I�ɩ��ٺ%t�������ŀ�ɱY�ЄY�����d'iMb�����N��Exk;N��!�������w�~=�"[{�h���5�,�H;d�,��rS��������/&�ٔ*��N2���#�F�e7���?QYs]d������G	��LM�Z���6�֓ԇJ���ڨ�Y���i�5� �^4�9}y�?�&��D�T���c����V��;��nU)�M�g����"�� j�@�5&|�+P4Yi�a.޾�qkx��(��o{���7�-�Qѫ�sG��1t*�
���^:���wT���VP��g������N�r����`����چ���T�@�Y ��������Ħ61ћH������Go#Ã-�z��ST��l&0���ӿ�M�6Vm���HsR?��j�3��M��Xr��[$F�܅R~�S�B�J���ϲ-���皰w y�&��\C�=$c����˄�������M��*�[���uE����D�0�^n<e"��ˎ$�63�������K���q��I�/2%��q�p�B�2K����&�������P�������߬NmaN֢񼟟�.\Ъ=����*�t!�ft.:�&���]OIZ�~]Jٸ�v~'�����Ɓ���� ڵ ��h��|>X��oQ�w�g&⛀pTʭ����g1p�<��lbʒUc2a��/�ސ&�m��B_��!�����l��S�q5K�Rǳ��8lFG�����~=�Td���V�!���C�N4:��k��*_�󋙖�9�ޚe�?�����4b�?�S�d��d�7���98��u�\�U��u�xW6�p�}.�7�m���#և�̄�p��;�S_6�Dǎ��*�@�����P����6[�i�-��2
u~%���7T��wEi%����!���)���lFq���T�h�>��.63�#�7;����
qa����/z�����*r�a^�:���o�W a��a�����uW�ߢ(8�I�\�D�j�����ސ-vc�#V%����O���x�r��Z�=Ed��N�dn��
��5mZ���5���mP����J�fx������Ş�r��{5g���z��*\����J���<�|f��L�I{�ܭ�JF�do�c���D~�Q_������tMش�y��k
~P����c0����ͭ�I�-XpVf�S��a�TJ��Yx�>��X�0t�����$�y�$��B�������T'�TڿezJ��d/=AN�,�N(��IS�9&k._����m-	���\i��n�:�eÐQu�O*���[���T���vs-�͝�^�\U�ձ1vb���O8�+�w*r�-�e�L�������d�J!��ղZZ>�{���^[V?�/-��C��ra�l�P��|jpS%�70�]f�hP)(s+�#�|�a�8��3W\.ҮX�	�x�u��;>�უ	�����ɩ6RL��/��7�%P���x��#!G4��g>�N��Q=!�0�w�o�W4���~��W@�h����rc���E������@�n�ئ�Ţ�Nۯ5�Z�2*"'�bw��I��CU��Y������g����B`����9jN�oeO>�*#����Y��hF0
f;��.�}���ي������ω�
���\�0�+\�T�?Id��P|��^o[!��|:+��uHa���C���:�����3��̛6֦�5[�ؗ��Nn|m��&�L�H��i^�l&���^��9qE�>�������8ೋ䀊I�@�bhG��P�m�=��e����H�Rz�(F����A<��>�hc�0䱜�B{W�H'Js���~�q:�#V���?`�=�rtxG_�����E��G�����.�}g~��R��}�l�^�Z��S9x�"jB��?�d�ԉ �t4F�k�X���˄h@(OHO��Y��k����
r�aT�pw�}�!H�g�i	�S��+��4���Gz׋�Ǿ����ݧR= ��?hA�����)�S�oL��L���yr��Dl��Z�[�MIUªko�	��މ�;���1r�Q����v�&0)w�Ԥ,�_��]|�ã<�1NJs���rH��Bw���ёa�ΨϨ����l{�PB�A�~�T��V�C�>~=���e�X]S��#�&B�L���2a��%�U�� N���ѼS�.�a���d�j������J�NU@��u/҈8�Z�&X $e���7/�q�m!<�wdt~Q<�d+]3��,�ܫ�͇W�������I�~�A���X���BT&H�!tC���i8�s�k���f�Ϫ*�y�G�W�q�@+J��M-T[}�Cn~��Ļ<Iɑֻ��^��5���P���O������>�߻=��(zmh��Et�YmRj#O�����^�s��%��Nn9��q�v����|�:#=U>�ȵ]������m����Y�|٨�����O�0N.����FğN'�u�;�,�s:Y~&����1����爆��ľW�(�:���{�r��(
`R��f��~I5��9y��:o�m�7y.�-[����~�+���0(h��������=��{�א��u/o�e����o$�b�W�v�&�l��=E�B�#���N��ҩ�2[�w��PP�:�eC2W�,s#�о|�_תk��<g�z�_bB��EL)�S��+�n�ݲ^��|�yk�E���C[^�N�~�ͩa��n�^�\D9��c�#�<�,ӷ�b���H*�ǂm���7�u��Z�o�t%�P%(��������׊�*&��񕛎������h�jC�-1�=�1_�E�t��~��#Tn��p릅ֶ���;�[sїG4~�Ng��	K��K�Y��'�!��f�b�*�G�n*�۩�﷎�(N��O���/�6j�P��a��7µ���:0[����|�)��o���i(^$����wC�ZZ�t���q���3+D&�����,�+y-��5CЫ�VO��KdpH��k�
�
#���3����a{�� �b������f���M:b�+ٯ��?���+���c�	�,�V���Q
�KN�f>J�P1�
�% ^�}չŷ7QL�=R!����Bu������$d �
�}a`�<	���Ҹc2�Z�oz5�N"p�����C$�����%u�#�x��|D,��-�k��D�jr��s�6ni���n��*g�K����vη��ω߾�J�����c��ir,z�J
��Iyct>�/8ЉK�L�km�.��ѽU�l$<����GI�Up�;��aG�l>���+⩊���R�t��di�7����a{�2��yx�8�K�PìW�MTD�eV�B�p\|Y����7�;��\�W�rϣE���H8K�D5��������hy��"vE����f�J�/k:�V�{�p�1�2#m�l�<��Y-|E#f0�M�5�0��X���-��p������#���n�l��R*j�l���
JJJdBљv5Ya��Q���e��W�*p&�K����%�:f#��ϓ7��z,���������y�L��M�z��la�yA�o7~+��(7����<�]�ҦW&�N��[�8�u��>έ�<+�e\��U�����$Y��ч�).�")J�?X��U�p�N
����-���
�L�.,aV�D�i��Z�����t�r�o�����Pu�[�a��J��?wu�n���w��-[.���q����'.��^��������t�XŤJ��i�0�3�ю�}��ק�m�,މ����\�����P��o\ 4e[G_�����P��[��7���o��rE!���"a�V��7��^Zpe��M
��܏��{Յ�F@*wǋ�S���t>�F�U�����CifY�g`�Sҧ�}@BT��Ϝ�{�2)�e����YZ22��Z���D�a�� �2��i+��=��P�g�3#������:r7~p���W?��G�p-t
�:��pJk�b�+�5w%�߾�b�9_�xL�'1�)Ԝ�� �i��s����# �����;0���~�Ss>��6�Ѽ�d��4��VNY]KW�
�<����l�E+i��Xz�4�4@3�qyr���5n��FP���'�� ſ������b @ß��Ϧ��~��[� Yԍ.\�d��1����D[�s���Kˏ2�X˭sU��i[R:�@'&�C�T��z8mXj�ޗ��8������op�q)��6�{-�~�	����L�~P��Dh�:��??����~|��K�V	�yH@$��6s���Ԋ7�����L��t�&)�q%���	���	���n�2��5X�)k��z	����G�}\�p�jQ��ecg35LT)��奜�����R���݅�$N�vz���W@�o��뛰J9���?^jsU��etH!qDt�	���^��g(�D����{���.�\�����A%�7\�,���
K%��~=��P��s�猓7���FW�GO�J�s[2��|�n8�wm-e�ŋ����������V�?v³;���|��d�Η�S3���-acŪ����wW�&��[���<�ɺ$�����!��`���Rc��ݍ��_��3!��Si#� {� �ae�ں݇��o�@0��s�ږ�e��O׊-	S���|vmޓ�^�'�q�C�m}�wr��~���+��9wSl�0��{�~���y!^k�^�[3���n�9Cs��6�d*�ZLci��}��D��"�I}�6����s��E6;�!�y�Kw@�A ʧ&�YH��ܧ����ԁf5�b>��'����l��g��М� �i�r����'{�IV�5�T<��gv�r�vz���>�7��'�%�A��
`ρ�w����3�F�Sk.\�B}!�ۇ=��7�u��ײA��t�[w���#%6�~����\�������>�-�K$�{9�!3����;J+�ލ8`z\��P�A��=��@]ߞ��w���PM<G�{�Q��skKV��\��<ڪ�?�@�#LIt�7�ZU��Q��=۶G�UU{��dC���p9B�|�ê�{DT|*��{�V�m�O�Տ�▝Jl�%�Rv��i7̫k�:b�U�oЊ��K�"�"�F�i�Q�(����p}�����d���?�W�>������GZuv���6��'(�� M5�hy}%�_�sz��G#����� ������S&ϋ�I'lK��x��#�r� �m�o,�M&U�%��<����CQ��/Dm8�t׳�]ۤ-0�O
��B��O�-U�`��q���]W��8b!��*���g�U�t��>xuu�v�ݮ����i	źXv���b��=a���@��P��[�.7=������u-m��E��?}�^�_�ħ|�B ��%��YD ;��+����M��-�����ws2Y�A^N�A��I��Fvg�u�ԁ=�IENA�vt3�^H�T�]��!d�%OX+|`���
:,��
� M��8���ϻ��JF�T��о-��/�Noj�����hǠ(`�ר��y���r�rG ��\�����V͈��Ǥ�W ���}���a}Zկ�I�����x^�Om�mм�O�C���� ����>�t��s
Ρ՜�B�����vn�0Z�u��c)\��4��bnNK,�i��&�M����u.�t��C���X��d+�i�d�?1�;:���s����c�6y���'�t@$�j,,=���s�\r)Hη����+�5��=o����T�	��2C������K�Ϝ$N���!�ttL��NNI/`�W Z��c�����yk7ћ���ٷ+�Z����me3rq�I�c�d�ʰ���l!�bC+n������3�zH/��奥zϗV��~�s�:����\��U� �(U�\���r�$��i�qLPS9��$�SH���O��5Y���w��{���M{p�j��|M��\��1�0�3���c�,��ࢶ?
���HH�tK#)"-���4Cw� ! ���90tw7CH��1<��O����|8���^��;{���eT�f�ڔT��|�!�#�/���-g_��aJ��aQ��3x5)�z����#�sθHg�Z�S�9l���ǰ�b�l@�OKݑ���X�_<Z
?�P�P>ԙ@��m���w ��az\�9�ƀ���CW���ږ��=i�S�XYY��į�P��gS�y��D_�7"e�u�Lg�i�4���i}� l���h�U��g �V��Pu�����H�3Ø�����P.��yVII�2��'�{�WF7/����n��U1L\��le����A:3o��E�S���&�.&��h�$_��S�ß� ��=:j�PU���[#4q�\���	�l>	�]s�<bS�������ԭ�[C�r3���l�����j�C����3��+��[)���A��s�p��[��&�c%g���`-Ok��W���zU����l�$x}�KNv[��g����J����M<7J����T�5�e��p?�w�$˦��6��=�l�,Ń��z��3 ����=�����њ��
��?���f����eSk��]2u��i2IX5z�V��J�z�x��a�]�ͧ�b�J�jv+�#謝��T7���%ғ�
���ċ������8�A������y��_�8�N�mP̓��I���a��
�Q^�_o��^�p��/ĬF����uxd�ނ8�O�}�����<���?�9D���7�}?���e���k��2�C?1��h�$��m ���~ǝY�rxu����/%'@B���ܵi�*e�V�W�9�cmm�S:�ǕK�<�;�ﾭ��D�ʹ𩑳n��C�lv�B ,���0�y�pq�`�!�v�Ć��[6���i�1��6(��J�m8\����0yJw	�����s22�cQط�A�Jd�����e:����S�<CHV.T#-�!6�k8��'D�eq�1[�*i_U
2��Xl� ��]�/Ia8�G�Ĝ�-�my��߽�����;�q�E��8�/(��ThC:�-_g4K�eMO7tڟ n#�{u�%�d��숗!�*�QgJ��0���"4�^���A�A�3��a���f���_F���"��ԘGM��\j���{��d��+��Ѩ�"،_���Z���`޻������
8�n��n8��)��v�r��kb��׷i�I����-��jDt��怖��~��j�-"d=����FjF����<d��?C���1&��B�����k���r�R��N���ȵ����Շ}����ig�"T�#z�Om�VfJ&ߎߩLj���=��K�qu��ʒ�&���'���~��-U˦�9�M���ryP��a�`�<��{��%����3`�hw�Q��`Yv[��6"o
Tr�*���]wD��훡u:i	":Ҥ�3�_*�{#�K�������)L�"K�X�2�^��Nt�����Д~1bb:�sv�˕��-_K4m/���1V�ֈ��&H��|'�.x%K
O�tz�����d�,y��i�v��W.)Il����+0.�Z6x%��_ԋ����_d2b����Ɓi���ܰ�&���9��$��b����;>�p���N������s��4��I�j%hj��w�T�R-�9�C��\*EJm�ӯ�*��܍]f
��s�bz�G11�wƟ93XlvI)��C5{�\r��H���(��}!��
���lZ^�p�h�柿��OYi+d�#f�2b+�Й	��L���?�cB�SX C��ҏLŇ\c�UC$*�]m��G=�E���E26h/?Z��jy�d�W�S�+o���v��]���,�ֶ�]��Ĳ��7	���L|N�3�R2$��D�fi!M�eH�6�KyeۆI�Lϩ�M�����6\�_i.���=Z�-:� �vcb� ��w�� ��Mf@�B��Q�j�*{�	J�G-���-+o�,{�������?^�˧L��T �k�/6���������<F.���|����}"q�[��Y�k��xa�������s�t�#�0uK"�f@;*kģ����|X��"�[���I�Hn:Zc<�A2������v�`Un��'����jY��1Xc5	P�C�5�t��+�?f+VE��w���3k�p����"RY�)�U�����5����'6�mq�ѣ>|f
0���� l��U�	.Z������ȊJ2?���س���+�'W�*����V{�0�ܒ�\0��a9!��0�#n��^�<F��/}� ]<������5�ۖ�/�-J����R�A���z�u������'�OXy2� �l�P�3��t|g�}�Ʋ�##��D���/�)��`k-߻ˠ�
��CH/Ksǽ�:`��D��	*�}��KOR9�鯋�_X��N��Ǖ�a��XW�[�?k��#�!R����t)C��#��R9�0����*gܵ�p�o*�A�ھ�;��-����(�J��.nh��4�n����?�w��U���M��}���z$��2��Ֆꔨ���*�8����i�-�;�ϛ���9����+�e�-_ΐ���^������uXAC���~]S����Z赋Z&P�����#&�Mr��"�0�N*� ����rƙ��b8��,�w1ao�ⰽ���z�?lQ��Q1�݆�=�Z�`�J+rd��dAp��M�F6�����32�� ��Yu�@��6��KC��̓�9�YP�Ý�賂P+%b�a����{y-��#�ht3y�g�Ϭ�iо��Z۴�{\�����$_�,0p*<��$���2��;�Q�.iJ��`�A�ψ��͉�Ͱ���՘g������W!.Z��[�O�g��*�����~6�����<�`�0��*A��^��wZ�)5�қ�Sr���uN��-��d^%��<t���\�ǃL�wCBQ3^8HzCݏ���`��j��y����[8Ēֳ��Y-)^�����f��(�K�O2Y��LޅL�p_�>�N��hp��q�<;p���D�����]~��P����H~E�����IJ�"����@g\_��Ue�'ց&� �[�x���x���4�=z"E��)�u5�ߣ���Q��ϩ��b��,q,&*�?u��IY���� {��#�q�5v�Ե,ZM/��~���&��B��CxAr�<X{H��X�G� �	*0yQM�	���3�p�c�nɆ4I�ghu+`�m~Ay3ؔ������
�P��ȟ��r�f̎@�y챙Ts��l焆�1N�),n��^uW��~��>L��R��4����D)�U"Fu��MO���܋TуSf,�\S��2��R��X�:�����y��s��^����Sn���v�5��M-���LN��F=�@�kQ�"�/AO�U��i���쮎��ހ�q�ؐS�ʹo����xse�G��1����s��{]�}G��)��x�P3���n'u^�k�O�10�C8aa�v�5R{nFU:��x��d���ĮbMY�W�Ws^X�?@7��&w�[���n+�����<R6O������C�	��YKA���,&bV��&��XPd_�|���$HB3A�g.>�#��VE{��V�Ǎ�K�����Mx$���sKKu�"rѽjRl�~q�v;�#�u�*�r�Qk�A�5A�dV^�ZKӑ5��%������'GM�[s�P���Z!���V7�(����:wX�I�+������ɘD�k��AU%9J�
STl��P���]<㚨��������R����bW!���7��?8�<��p�0b�~UQ^gS���o+Ut�
ޔ��3�.���w��y�G���P����-nf�<�I�t=j�9����h>���}P$��^��t��m��f>�볂q*�(+�LI�p-�"��`�/��L�S��E����ذ��˴vv ��^S�f��jǞ�)^�wH���:*	eaVلs�t_�zsi>K�gp��'�MU����]����EӚ��rQqz�6���[L�l&��g�#jޗ��LS��2Ü�xh�t�t��c�����v�8C������䰯ߚn��q���g��wN���|�y�]�FoT�M�u���h��������#o.&c�q
����f~M����$i�|��aO���9������ly�sJ�8�حOٗ|-Gk�|�ue:����3���X5f��5��-���t��wl����&}.
���Q���ն��B5�O!�'��HV(����~��"��@_H���0o_��i[����������^�Lf���T����T��1]��L����q�{�A+���N����wX��;�D<c��!3'5A2��E}���j��UItK�X�I\�V�Z#1�$a�"$�rr���F��¸���8Y����|b/�<2�g��4K95W�jC'>.���?�XK_�|���6]ؿ�}O�[w��	u���)��]���t(z�C��ek���x\N�S�n˄v����,���6�'�~�nD�s��a��'��e���UR�C\�9W93��Rw�{��2���<@��ZZ2
���EhS�gӇ�� ��81NYI>�WN��zScS�'�����7���Q�"��^�B��`q	CW�$/��ֈ��k�!:z��P#�7������C�K4d��������ic��t�,;���I+Nڔ����a���W�S�K�s0J����B�;�g������Da?��S�kbuHu'���b���3 ��!!}�����k���Q&Javr¥/�4�=�jV�+KJ�S�f�T�cASn͜�/�9���î�Z�Eȝ�h�m��S���.Z�[l�����T�rIaɿ��w2I�^l�w���A���
�Żl�JQ&~'��W���+����]F��@�ip^��U�J�˩L����;��Bb9yU�FH��ɒl�������8/���u4����8?�u"~\[:��R#
�a0��[^���F�����A��yK�v�w��/�;	�[1`���߬�L=�r������9ߊ^��[�p�Q�w�/�C_��2aO�O����A��)��F�A"���:����(�~������?��">��׻Ģ�U�d���;�?JG�O6���f^�г��4����|D�|"��aP8�x8ļ���%���:�i�t��XM�B��i{r�G�WW�n[�E�O���V.N]ø�L[c?�˜,p� 	Q�Z>�w�Z6ӓ/�(Ó�z�23x����ZP�B~���Yl�k�����;y�8�-���o��]u�#���ҏ����<7��T��I��T�!t��h���c;�~�[�w_���BU~<S|)�h�,�h��ӿs"n�/�}~p���q=-M��E�c+ʲ��F�i�Gw/����tU.�v�Rٖw��t-�c�\�^r�'���ŏw���NW�l��x��S��Ufh���&�Y������8�9�h/v!?}�z*K0����J�K[��r������0��:�﷤ɒ��;b�WE��O*{H-�]�e6�D��ءQ���Q�����f7���q��5YV�=X�c�Z��@�eEE��~l�!x�t����H0��;m�{)��A�sǶ�[�xBm�5-~�m�o�rR����u�=
[P�}�����;
1�I���_!�ꉦZ�YDG=M���(�����J��������o����u-�\<�eu��s���\�ܮ�oA��Nn�"�(Dޕ-4���6mZ�.1���N^G��*�O�1���u�W��t�X����'�<u=}I����́�Ƒ�i�7�5`�U��r&#;���L5ܯ��Ez3*W)T�5�I�ړ/e PуT�i��}�o@�`�/F}�8p���2�����EE���;���ƤZ/�}��Y����B�J?�U������6��0Z��Z�s(�&���U}��?v[��QV�@��Di67�gVN��ZK�/�m��"�r��Zd��+�bR���(⃩g Sjr� X���§7�]�|}8DjkSv�{FV&e�k����q��Hf@�?܅�ɐ*(Q����9@�
�n�#f��T����W��)aT18�̢N<v��SS��=���#�W��߻������/_kC c#��F��>!�~�R�^摸S�6��N�=����®`!�\�
����1wy�[[+�H�n͆ќ�B2��1�#4�d?�8} {�ɝ*�'���,(�7��χ����{�RH�����s�Y ,3/,�����×�)]��T]�x?����!4��JV4��3@�3~u2M�:�c{��L��IT'�����?_A]*p���`��:F��<����w^m���`�.F����'U�~S݈����+W�>� 7J���d��+��NZ�_'�πK`2����]xF��Zʋ����>�����[M���b�K�L9���N���B!��u��c��d`�}ǒ��iu�����f�G�c�z�(�+B�{Ww4�|Ck�ӈ~�(��Id��I)�2�N�6�[	��&P�~�vL��E��2^�,4�ѡ�U;�D_��§'�7���yVn+���S@�I�km���/��"^��MπM��0�����"�m�5������Q�Ydb�l+����8�)�.g�'<�7~�w����ד��ì& �����C�`���L�C�S�x��^G��k<V�Q�yV�OTe��׎�']���:վڱ~Y�*�;��V���|�#gZ�t4�����3k�[(j�ѫi[	���HCw��	q!pU)┣�BT+�9����L\a/U���*�-�)��4"\ <?Xō�']$�j�V�tm[j�/���?9���cf�O�vӐ$�^ڐM�p!� �挅�gO☠���z[>�]��򧋀��T���Q�]�oj)[��ᥰ��C����	j�8�|�UIu�b ������O��+O'D�E�&~��z�O��S'�n����>p�>I�0�E�O*T�����h���z��[#��Te��tP`Z®��5�� P�.=v��-��Պ",���)�ҵSOa�G&�w���Jet��_���5˅�ٰ��PWՐ'�P"4�����So��H0G/��paR���[M�2��c^���ՠ���X�U_^D�y��J�~LE�-��.����B���&��1�+�|&k|���%6�@�����|X3���[�0���'f�5[̅���ļ�Y��G?���� � ��M�0�\\S�(
�mz��`��C�z�D'_��6w�Ee�5����r�+[����0J���%�Z\B���]��88?H�d���i������B���85R�I�K#�=z��)0�3`��ߑ\(l��|�`� ���+	,����z��f�ྉ�?�Q�]�r�2U����J/Ǒ_�/�h�ӨV�=����#��ٲ��C�z�JsQs%nT����h�?����tH``�c�+�g��j�ɪ���(����ľ��8��q�x���������E�b���'o���y����1k��A]pi�~/�%��q��g]c�.�#ˉ�Y�P������{Fx�g�sm}��[ɟ_`�v����$��1�R��p�1��L�w���
X"�izv/�&i��Hy��b�=6M��<ܳ����-$�m�I�M�Y�K��^;gg�K�䠊���L���t
��!b��X�����KoBi ����!e��0>SI/�&�|΄S�I���#�V*mv�c��NZ꥓҇n�P�!O�_���8�k$�"�7M���
@�$8V�e���i��X�{,����]2F���e����}��؍��{l�B$�P=����څy�7���i%��Lԅ�I�a,�DI��Y��?��z���h�稿 ,֬��zI�&���'n�Y�I�guytlXI�k��ι��C4�sd�͢�M9��m�Յ���'!�ƃٺ)����z�dÓH�U"�b��٧l�F�a.�+Ბ��z2}k���4��F��n������b���4�,M�$jXk�_^_f)��u_�	YPQ떜�b����zx���ޝh[�
%K�c��s$
$�*��f1��֑&�~���"i�������3%�٪�N��r
NYW���7�\�G6���80[y��%7��.V�	�t1a�a#��1M�%&ț^Qo�)�:���{o��ؙ).}6�!���4��E�oq/��B�|	N|IB�.x�ņ����g=���X�o����"m�x�.D�X4��RlcO����2eZXXQT8��/<���@��:�T�L�i���L�):暛xJܭ8��g3���(sN@b=��dg�%Ì?2IC�	)�̎/hK��pC����	&��>�#�%�?�*e�\��-��Az�vo���G��Ɛ�=���8q�$wr����]�F��t�����q[�j��6���D�P?�R�i�ζ�a�����ֈ�C�ʓ���2[�gs�ܣ�ʷ+-K��6��Ou(�e��������en��������9l�z�q�	h��K���͡��{��)�[��Aa�m?Ʌ�/����s�!��2ʭ�H����']G/Why�:9~��6�z9�x"�%����p�m�w�i�!�����.ޢ�~i5��K�,�N>]J_�A����C���F�ׇ=��`[(�����x�iz��v�~������y���d��g���7ٶe`9c�a��TW���w6�T�ن��D�ZGI��fگ�"��͕<����I���C�n�zv��KT��[�'��+Z�n㋛�b^>��\li��IS�X�Bc�t����g�Ta-oY�n���X֧��e�
�g���#�;	m�ms1��n������|%�:�b��M\Σ-kB��`�ث�/�;!�g�4�_�<d��agd��N���e �i.Aee�������l>t�������֑��?�*�k��{�|�ڹS������#a�Lv�U?�|u6�1�Q2�������qeK.���U&��.'�BB�_[�|�b��u�	�a̞�Y���z)��>=��z`���VE��������(od�s	O~������͹�\Cy6��4.ׂr^���j�͎HƵD����d�˰d,q#rJe.��p�/�����[ߚ�ݙ�e��c��W.�H����5?"9�){tԃ����v�M���q)��~�J
�q�V���+�GQ�+l��м�t�`���Tt)7�n�A%��FNJ	m~���e8�(��;cE��낥�������	���H�?s�Q����������$ש�3��K+�6ɘD[M���e1�J���F"�5��O���A�[48ה�Px�<�y��>�H{�=��O�ி�~c�~�sGڏ��>�c����4�ƭϾh���7,�:A��m���U�|��Ÿn�/}ّ.������C�Iu�ɢ>�����_ֻp���[�&����D˞��⤫�e��A�W�b+��&/�US�h�h<O3��|���L��n �xw�k>�})�����JGO�0�(G"!�L�����"�I�n���72-��5jc��֠d�4OO~+PG�#F��M�+���� ��Y[|����Wt�=[������$d����VE~��|���{����!��PB?0��D���f��/��|���O&�)Z�l� !��W�-�лe:֢1]�H7�w�q<� g�?Q�7F����lK��G�d�X��J���m�D��8{�HjQ���!]lI���|`&>�C��SN	�5�Y����H<\�s�U�|�1��%�����4V�/�É0�O���fo���{���:(��
��� �6��p��\J�Ex�>���qH�/:{�=��mC,�h�Z�7����O����9dWemu�/=C� �CQg�"HY�\_��UF%1�~� �ˋ_?U0�x�-Pzص�R�����km�����USL�B�����{@����~/8>1���gO2���Gl�}�DFm���������V��}1��F";})ˇ6������|�tpy<�=�(D쾺�Ǳп�gc�f}r#]���ֈ����N�彲1�"�>l�X�G�A���b�}����v1��!��l����>�Q�<M��Ϩ��y]_����స���AOzE�.���~���(��;p�P�?�$!�w�Y���?����Y���}ǚ�a\�����o^ذb�����șBᩀ:�3���������促yQ��J.�!�y!�����R��z�{#�]&�=�=S���) -�my������I=c��1�(���-���!�.Q��7�krLo� :��hiZZ%/����eux�RM*e�LY�P��M�h���������%$���6��>��C!�{�yä@�Bߎ���e�{9N�(/4��[A?Z=@E������˷��1j99M�@�{G�
٠�S
��_=b?�n���6f��䉈��;b��`�"�&Dl�E�&��MV����/�
̆���0�"C਱b �_�����mMGm���Q�4p�426�pa���)+I|o�������{&�
��p���[�ճu[5��J��J&`����.Q\[\֟�1˳�^Ҋ!�p�0�`�\�`U��t�'��V��}�`PLN]�H�[�E"���Γ�&R�Կ(Y0Z��3P��j3����J��eGI���?���^��bZ,��W�;��j��34g���P�y�J%�&�̷�7��D)̍�uB �Lu�VoI�������(y^�M�.�M�X�R���:�X/�G��T���}�r���lc��v�w�f�o���׸'q%;�;�|�ުg�몡�T��VE:�mL�֋5m�tS��W�����Ԯ���E��j򋔫��ak�d�:�"tn?0�*< 1(����:ʼ.�ERW<�uH�G����W`~�K���go�����ݛh� {�V��Z��悳����T���wt�N�S?�/���L\��ec��X3��Cr��B�M�l�*�:�W��Q�_]��WG�5��y�f���U7@�T��"�
�l�m����Ŀ� ��[�Ky�P�n���d���p>*��_�l�QUTB��k�������+�V��?�0�=��
��6�,��e#�4E�j�d����;�]�V��!fe��j�Rِ�ods-�x9�� `�i��F�(��dr������R����1)��=2}R�F&!�".�$;(�K��΋�TM
!���I�M���u��L��O�}��~z���:N ��Q!@�Um��Dj��}-~0x,��q�������$`h�$�k�p*~�����<5���[r.|�TΪR�^�ĳn����O��]��E����W��Bb�w��/t6?�X	�5k�i��<PVk����;y�K����[�+���d�c�[�������9��1��c�],����s�t?޵�:�,`�F ��������X�d�9kŠ٣���x���D����=��E�����a[< *��xE��M���Lʴ�ݖ�>G5� m}k�
=���l����7�u^�N?ۏ K�_H�t�����M�:ר��U|�A9\��U 	�a�v ET�	��s^���gb`\�-syY�con������R�cԋ���a�a,�$�f1дC"�"�X�[%L���O���I����� ��tk/����$������#�!%�::\��H?�u��k��ua�+KK��?<�������rg|�˕���.�����x��̜���߮�=j�,�T(�5nE���!�Ub���'Qݐ�FE���d,��#���yq��a
\���p˳��d�'�,�F,VS��n���������w�uM�ު�D~x���
���wZ4�q�gM_zХ��k�����^hV�?,̳H�qݵ�{l/�Q���+�g����ǩ꘏����>\<e�P�]���4v_��om�k��-%4\�u�yk|��VW�6�%��ŞU���a�W�5O�j9$Z�u���t�IfE^�V!��j|`@W�5���ef�h%��.1��y6����U��*u�⧇t���F�7���^b�H���N6���"7 �w���Y�7��-���Ԙ������9G����Ucw��Mb�B��7� ��ۿ�/b���6����{y#����V��>al4�Dm�<��&�� ��B�j��Zl�])��W#�9�[�+>�^6w��D���r{�}����B�rD�FVTN����B�ଆ�Ș���U>W��Y{%�����Df��~ #E�g�2��N����3����,�� ��#T�)3�`=�n�]Բ�s�#|�u�靍��:Ud�ې����L��(+�i�x��x��T��_��?�����m�FK<���n!ۄf�Ͱ,�����?�K!NWj���J'��q�+�HD(}s��}���u�asD�;/�;�XP4���C��VOƓ��2�=Z�����az������>.�0��`X���Q��#|�^��q��v'�26厶�<Ԓ�!�YM+P�sq{joù�3L����O�A���\����J\�Uy�oU'Uww[CJ�4:�����iw��҅�q�?�O��K^���嬢���-���mK�����Xi��X��\����~�	��5�z/�1K(�$+��nCo���c�k�E�\Y�MŪį��{[���B.�+[ia��~��U&�#NƁ������� ?m�'�:i�K�4��O����A���=2�� v�
gc�[� v �+�.z��nM� �4��:7�S��4�U��^��L�Ri3�����F�����k�m4E!�%/T�!�\Tr�cH�7��PIW8|1hhhj׃F��o����KO�U4cZ7��O��T7�4���.6�ڵ��K3#N´8Z�s�dVˀ�֙O^(��p�a��qy���M�a=k�]:;ɩc�ձ;��\����4��?7�Po'�S�{�x�;���_���#pڷ�!�I�p����8�u�5��~mlw[h�s�M����|;�&�u�Do�9����SA�+�HH�&��ɱ����S�F�z99�����-��1�O����6�$��Bn�:uH�����1{�CY��1�]	��T���P���k�@�?HZ�{Xq3���Y���clҠ��m��艑�9��u��E����鬯��`�l���,� ���z���R @ჱʸ�I@����d�Y��V��@h��u��w �s�&��G�t�p��l����I�/ �a�@*�ȑ�����Ga%|-��+O�q����;2�!�}Y��_q�%�n��Oq�y��㬗������Ɋ&��݂�i]�?	�;>�d� ��g��f��q��U=o����*��Or���UH�W�BwQFc*{nQ+�7s =˦��
}{���^���W���G���\�"O5�(�����(J��?1��vi��ǌ[�?�;i%�0xDN��=)���=�˜�`sY�����#�J����͘����������e���zǞ�'�"�����h��EX����A��T�ҥF?��ok���R�!�v����t5,o�A�����k)Ǌw)(���6��(�F6a��S�%��E
��>���'JE{E�R@��鰬.^��nR9:��V�/T^��u�O5�OKr�{�ʡ� �|�N�e�Ӽ��?w���#�7ҕ�Ӧ�T�(�v�ߜ��V�b5�_����q��g�/��Eű�Ga��O"U������M�����4A�@����Axܒضm�W#���"�#�������C�����Fn��`T1�is�T$���_�w�P�o΄l@�����q��b��]?|t�o���%K:��1d��Q��jk�^�+V�c�i8�u眨p�5��O;��0���OSh���^��ԭ��yI�q�J�#�S<0ӡ��Uʐ��Z�t������{�$�RI�����$�ֽ��j�'HC�N2���)?�u�$#�B?�_�F+�-&���M�s���L�Ď[�=�q�?*6�2g����D��t�-��eB	��O޸.4�π�I��B����sH�EeE�����QS��J݇�?�ta^G�oVR~��$1��C��"o�S���]O'�"\�p��6�������r�V�+k�gyM����]�L=ǔ���]s������:�3:Cfuߍ��pO��g���>�F����r��J���*�([C(�FnR�3�כ��\Tb�����}oTn�������z8Y��ݾ��Z5 ���.���AD���DP)!�=R0�\���$BL�NY<���Cs�>��1h��o38(��\Ij��i�����t�a[}X_�bR�<�+�O���lb�Q�YKO�(�I�G�;�x���Ow�F<A�Ӝ忇o�z�h�hb��+�-i��8�n�mE�P�1�W��h��<�|Ps^��N��l���QV�MI�Uʒ����ߕ�dC��>��V�dg��O�����;f�����Cf�,��
� ��g��g@b�=b5x����0x�0o`��O$�ޫl��MIBZ�#��������7g���vQ��g�&N�W��vi���!���ť�I���	T<�$���1kݼ>Y�_^�����5_����5�6����m7��� D˦��:�?�����cV��U1�r�UClJ��N���M�;ON�bc��u!W{\d����o;�����FGO��,\y�����'�T.*_p	:��;󽳺mvW�ckâ&��EC���w�r�C��h�XW�����F)K��LC�bJ��hc\�f����".�ЪJϩ܀�Zl�({厎����|֑��S��^�dU��=?W��а˘��o���i�!���o��!*>�<w����w,��[���tE{#���˞�h�[��N��㽅���7�VV���lfh��� ��db�x��xNT�ǿ.�`�0Z��J�MZ�����]/?-������У�����9��  �����R����>��-�%p�'������uO[���I2vb&����W*H$-+�܈GN&J��T�����p;_Z��=�g��&�e���xǑ�w&��$l���"�u��֒�(TY���aQ+�T�Q�1C� "����+~-n�l��
��[����ڐr2�v`-UƵhշ�#&��[���"r�3'C�'ѫ�����KkdƇD�cπz�+�����?'�N���~������|{�웖�A��,i�ޜ��=�W�~�W9@�BbK����b���/{W��qtss��5��(_2�ոW�y����b/��ڍ��RW��G���R�i=����XG���7���w�o±5�8N������W۳,��
����w��g@��M��iu�3�U}�]�e᤹��[<4�f�J�C���T��Z~��~F%��DS �p�pk��Q�,��>�B����5q�%�vJ-�� ������r�aD�U�4�߱�P/�$��UC�2K�Z����O��D�N��{��UV���v+��x�O�:��|��Y��Eך�<Wƞ��׊���B�Lھ��9��?~W�B,��Lg�� ����ǂeEf�1F )�N"�m����u���rg#=�A�/dN�"�i7��l�/wN�,;�p�F4@��K�x-����pJ?�4�'�wQnl�џ��nm2�J���4�j��c��)�[~t#���I
Фn��g��HH���A�g�]�䐑�T�k����R�?!�wqI�;N>;l�d���7-N������v�c0�y��gRv�\�go����J#r#����8��Ι��0j�_�V��z+��K��1����Ɔ�ހ"ۦ��49u����Ǐ���<d�L��r�¿u�Z����Ҳ�Ϭ���<g�>��BZi���Ώ��?�SOt����3+��.j\(\L�ܙD�^��#��a)|��!?����|uJ�h�Pd�]s3XO�~!ۍ2>��/*�`�یXi��:Z����r���,n)�y7�5,V^^~�8�$QM�dTD�D��f=���`�J�s�؀�_YU��ar�ȹH�_Ӯ͈���))���K��s(S ����?T�T����#��֔G^�߬Qs�
��۾
��k/~W�{��;��4�]YӠ����.�(3f�{=ThX�����Rv�-��a�nH���:����So';�n��Ϲ'ᛙ��˷����a5�fR�zM��g���O�`K@-*;��}�:_'Х�E���w�8/����K��^�|��=[߸஫�:�ik���?̽UW\��x����Np�����и[w���݂�;�ҍK#�~�3��{��u����F��Ӽq��w�P�o�G9p�l5����{߲��;����\��˰�0(^� �ޕ��vO�f�ZS@� 3_��[҄�J�R���G��|�� $^E�*)�����S%��+���w�P_�`����:�DEv�pb;�<�'(���ru؝����R����?�Ȋ!�KZx��4enm5x��i}e2o=����6T �O�/2��~��y�>���j8V�j�P/���R��_7������'}����^��*�{�����H�\~W�J]^~d٪�O�jme�����B%?���(Z��X�w����P�-�w�h�hz9+711ݭH���Pу%���w��[�{��5(�?����j$��^����������p�{�Agp����ų3n[�8WzG��������c�O+�����ڴ�)�#���'���"�e�m�o��66~Jb
�d*�ٺ3�d(��`[�Ӕ��L�C�<0��� �Q����TA�±I�GRI6n�i���	��f�Pn�2n�$�Se?RK�Rs��K�M�s�FBQ>R�$ɳ�s,��h�<c�$O�#��Cs6����i����E�A�U�[rLh~L�����bץM�[�y!�şP�e9f�[��i��4�h�EA؊24�}�d�\���[��,d�'Y{e�;���[�f4
c�?���䨞CW��Á�=&Ui=g���i�9�7h���}�d�SW��P�Z�yK�L~i���qs�����D"�OT�a�2y�R̗�������@�n8}�w�a���w��^3�i`�j����Fl;e^6��Z}ᛪ*�g~���|4������1eO�����*Q�{{�6�YbVs�3;Z��_�l)]j2t\��+�z�=��ů����j���v��<�4�K�.��f]hg�쵉ܫ�q�f�ņ]]��i<iÕq��&l"Z37ZN
g���~��"/B�茕����31�����ͬ`!�
�x҈3%\�x���X��F����!x��?[%��	�Mˆ|��3���+��}.1���:M÷\ԓ7,���2�L`���;[5L������z��|0�K{`�ߘ�hdɕ�J;�뿧]߫-��	��>��V�UN����A=����ڳ���蛴)������p��D����y	������g]�`�qR��*M����!�����Գ��Av���J���
��t�sÛ2H�!��V4��)�l�X؆Trh0�ۀ�R�"Kyx�_�H�Hs�c��[V�G>2W��(�Ȉ0iP��YajJH3(�l�0@D;���d�G�����l+��j��/�2�wyv�A���oy�z`�ؿB�Av��!0�w��5�Ը�FU����uO����b�G9d�U�;�J�i�m�.	�����"	��qo�����mW���tZ�Dt��\:V8��wN]puW/�y0��#���\=C�Lؾ���\���[]gvp����4y�e:�Ɣ|�!ʤ��I��*Ք�Q��H|��ےw����7j�Y��r�MK�q/Q��TL=�xDj��n,��ϖ6	�Pby�L��3���y�.ߎx���l �����8#��9�DO��J<2��ඓ�9܁��>�pY������$fa�ϱ��FL�{Ȧ{���G�t�>e��[
J� h�/��	�1��h��_����;/��3�	H�cmު�RMQYO�cT})�����~��C���⟑��굥����-���}�t��?���q* �}l���4p~���(bﯺ�cz�H��yZ��5���LM��KW�5L��Њ��f�`�����3J	��_ĥ�Z?)}#繚{�^�U'����@�ӹH>�|1�����B����Q�rmà�S�^$ٽv
Q�����/$ׅ�?$�~j�����¶@�v�� ۿ?&9��d�������+{]��F4k���c q8EB�╟����kݻ�<���@b��eD�U�0Y]S �3�b�3'��?�����=>ݱ.Z�U��Sq�����L��#�8�h�%xi���,D��a����a�WᎨ\��*�I�NŇ��Ҷ@���	'��y|�����(�%�o&?�NHZ�^���9Εoy7l���F*�"��&�'��J������U�$��tg�x�^������Jl����î��F��y6�L��~���*�d��:=
�8�tL��ԅe�xY�����8,����t�;��vDT~��X�K9(l����+�d"t�7t�?e�Z��~�\�B�y1s�i�6x��j�Jh˷l��=g���A\�I�TBs'��yI}�y����7m�;�`|�� �eJ6S֪��w�8��p���I���I�����V��8�k��;y� S��ax�:[��j����MMi�5;�/��m/gϐ?uٮ��+��KVU,�	H<ns�57�SxMW؇��������J��Dva2����&�j��Bd@P+d���0��@1�����{��)G�D��jo�;��"%;�gZk�ފ5��sF崭��P���Q�P��I[o\m����d�3�Ϋ�+lEH�T�"�Ĭq��S�Q�sG|� ��� a�bLk%Z|Lv���;`P��7�ی/Dduz�aq j}XK�g�]6x��\Տ겖6�=�ŷ4���[��cCn77�z��ꗹhՓ�ҙ���<PE��3��2ڍ{,{�-�'#�h�W��Q�%X;lЏQ�ǫ�����''j>����f��6����@^��>��n3�}��r��.�V�,�� 9�(Qsԭ[k����]��l���,I�5OQ%#�r>���Qh�FceQ"��zl��%�{`py����>��j	�]�$T�~�Li���Pe*{ΥFGW�."��!%�oEy��63���Q�|ag���D�m��`�ky4/�#��*�E�@�n8VuG�Jp	������Oy9�o&��uZ�0��:$7�<=;�2����Q�d�,�J�i�}0g�lK@��t`lDĖ�3�M.����h�P7�ʖRE��눠Ԋ
U�?i��9�~<_��7�ϴ6�9���'�Ne������r��8�n�� �>��u�J��~���M�4ՎCޮ��#b.�h�]Q����Z��%'�>�DW��͢v�7�*�M¿.�u��x(�������u�?�=��p8xGik������n�N~վS ��x>̖�x�Kji��������.t=�1��}=¢�.��X;���������Υ0����kk,�% �?�b�?J�x|�����]�����q�+����A	���CiC��U,X�E���w�h��q��S�g��$��wK�\kc�6`���Q3kX+������(�R�Ӥ��"�@��ʙBWQ��_�g��>���㙿�9ň�p�����D��܇��(j��^�p�p2�h�y�7,�>�N�p,6t2��`�ي�?����t��}�o`�A��p�0]�ƅ�����x�9�ʼ8��*N�t�;�QY�D�:ԧ}s���rj�9Ayt�e�����x㕺�:h{���0��Τ���2�J���֬�<fk�I��9���!�v�3�34H���_�JY��7���/���ee�Ԓ�4�����U��\B�\+#�/�� #���p��?M8Ғ^��j�5��w,}s���D#I��������MQ�ko�烬K�#֒Ԝ��Q��p�Z��-��A=��ȴ�,5��u9��v*~U�a_�SY�r��ٙc�qi� ��)GP�g���FPjX!�yv�W�KB����BѸ�u���ņ��A:�t�u[at`5��#3>�А����ҒH�����~�T)�*Ί!��<�J�.]*�9d,��R���ʿ
���d,�ӕQ��j�m��s�&��5�iJH�0	��)����Z���USA�=��FK�n�Z��aX�#��"������(
h��F̈E)�؋SK[����qzz\�hR����UC|<�>�_Zem���;�z]P�����aqI^��@/�#|�]���*�i}71ml���+�2��X9S�S�/n��9��*������9����O��iNƜ6�xG�C���F����=�>B�dhU�����b���'=B��]�@0s���� [)h�/�������g_p�j�e\����&:*��������z�P^�����4���Ap�ۮ���������(N��pޏ�.����L��,�Li�	�5-7���C�����;��nb�4����l�6q��D�����x����`���WZ�tO�ϔ�xA�(Mg�
ҋ���Wo/	S��Ǩ�;�ԝN�M���Ҽ(?���+ D����ş"�̟�j�����k�xZ^�(� 8{�,�|�WօG֧M�Q"����`ǵ}F��Mh�Ĥ4�Eד�eF�u���&�]cd4�����w�/�ubv�Uj������\l��F���5
8���6R�Х:�ۏ���bi��Ó�;�:+�t��h33�>�@��_���j��I���Y�=h��(��@��Jj
h��y��̴���5Ǜ��6�?*���=��0�h@��4����ȭ"X���a4�6�ژҚ?�J�^�Ԯ~$���)Ύ�N r�a���$��N��%�ˉ�.�t)+�H�a���$��/m���j���~��~���͜OP t�5�6p���k'P�������X���s��8�e�d����4=�TS�}��8����,1��\���{s|v�P:��Z�*b�T&pgt��]��g� �J7�f�([Q!E���muQ8��/@�٪�[[TG�;?-i�k?�zDC��$���C���uvb���ɥ���{r���E��qʫ�)�ĺ�2�$!�Z��U�Mҏ��{��L�
�N@3��\A]��� |�>��k�9���j(8(�F�m�b;���µ{]��o)hu�"�O%�kQ����>�M�����o��b���Ҍ7U�Ws'c6$��1l��Z���~��1�=�
կ�L���������M#�J��Ƈ<�Q�faR��@'$��+����Y��/w�e
�{��b����[���~��x�S�iOQ�Z�w����O
�\�"������..:���8:z�)c
z�\�'	�w+RJ<�Wc\�+ecj%���3:�$��[���Mb"n*Zs/̠Z^j�@pb;gN�નY�o��&�@U̅��Y��^����ߪ�|U�1eU�X|�CWVt��El��<E�j�,L-�F��^��?$b��H�G�R;���\ki��h�J�v��`�q�����r��b�Eq5�h���&�.�e������|�
��<�$7K���D/P�ρ��z^jXc��� �qqT-C��\5lq����YW
M���u���u
v���U��]�u1�U1m�+*:Rfj�:t���e���"
�����ST���(�f�l�ԧT�i0�U��*t�(4}��!D��Ul�ҧcd}�K�ﶒɬ��	b'�_���K���;}�{ϖ
/�	,��s�=��6��.NG�S�d9q�=~�I�5���Q��!n�7��A��l6l�+���tXwq��Q��4����@A˯�ޔYS�<D�K�����qG�&�Nc2��"�l�ܱ�����f�+�,Q�����7bs_���F���L&$�s+G髙�ҷ���w�s�K@t��\,N�O��#Z�-f7�q�]]�+2�÷��ƣ<wxW�n�ls
����>���5_3�	-O{}���tg�`��_��Rs1m9P��'z1-$�V���5Ď�����X�}D�5�H�*"��. ����;ckf���bn��Q޲|�V}��2
6V��D�\M#kh�?���^zQKkIq0�J�0 �-UjS~�P��E��>��j���<���DeT�+�W!�n��'mGV<��=כ�ڨ�� ���䩲q-��WSd��p�s^�!��kp�r�A]�_j.�"╟_'����,��nc�g8�o�^�C�3�֡��3X��i�Ϋ�[�q�����#G_Rjp	Z�x��6kGg����(f�D��Pr+�M_�V�s9��po�o*PwT֢�o
	����}�@s���2�N��2fC���61UcB#̴�h$��&��Bks�G�k0k���*�\�FJuo�3�7�h�Ap[uMp��x�z8{�^lP�!�=Dp��F����:�|f/�6�S�����m������oF*��-m�r����Z���\�T��M�_��E׷���r��3�A�NIj1�-CqY#L���X��4�$�d���b����^�v��K&��6�~�#��ӎ�p/a�V�Մ����'��p mv��K��ͥ늖`��;�%�Nq7�V�?��kYU��AH,oYڒ�Ud�[)����y&���7��d�f�֔�w�X�M�"A����7; �)跂���g��_VOA������}%*?�G�H��y6-nJA��F�Y�,5Q��	}+���Z��%S����ͩ�;M�U]�jg-�CJ�SdF�͹{�a�vG����V�\�����q_��IWMP������M�d"�|�YW���K��P7lx���i�g���ۻ��U��Ӈ{G��T��i���~&~NΫ��⺊N������=�ixC����<@�7��&]���A�i���Q}���\ڵ�Z5�����6"Oc�;�AT��bJvr�N�3�-�L൅'}��ǃ��s��֫s�f��T�O�鶏1��U� pP�bLQ�|y�����j�m)�3z�,rW�i�Q��3H��<|�V�s�<�ʾ���$nއ���tB���Ԭ���y[5$gF������~ECzIUr\<��e��H2�s����u����\�i�N�@��|�����eJ�`�2[��K�f�Y~<ǐ=�tԶ6`�pj�Ĝ2|��(��Q�ˋ�l;4y�;�q�Net����O�]{`^�f=-
,Ɛ��}wc��(��/7����̮r�#�/��Ԋ�����C���L	� �>V7+˓�)
�i6��Ӫ�e�������G��ψi<w#X�(��kmJMLm"{�m����⿰&#��a��� #��c���`�k�i�".>�Oc-�|���J��'����?M�Y�Qm(���V��]���W+�������2��o)���f�M���Gȥq��s)�[��p:����Y�B�;@�`W]!�)'�Ms=˝�>\���ofQڲ��YA#i�6佊��5�<If���5�-{�QO�ҩ*	�|yv�=���~�|�/��z��"��-��i-D�>&��Y��F�Zo�m�,��-<��'*�3�(JgI�h���9sH�d�q�$/�����Lo/��4�s����3�D���"���]�ezǛ���J��j-�̛�"�5'?	RE��o
�	�PE9ײW�	�p����E�[���i�:+��!.'�[Ģ�]%��{>!���ϙ?�0S'��pů~&r��%�4�dȗ��-����$8��>~���4z���6Q}�����4�;uj������L�v�V樈�WC0LpKt�+҂���Z���鹾��Mz77��<I��g��Y~4.|׼��xd��D��=��IUy݅`S�5�/��
�d����A�2�6�4�6	��nE[X���+��~�z(f�86�-�2ZO+��#��fA9E�\>�����%�ğp��ϰMW���8U���+����yC�&U�ߒ�#���ЎQǟ�yq:1!i�)��m�@^r�t�;�{F���J���y�*g��<2��?/�t��#���Z0-|����;`E�e��*����b���˙4N.D`G��y�w��?�Ҳ�g�� �F�n���&�x�Ll΃т��D���:�5� (mf�<��`qhi��K��HpH^?�v�Ύx�5�)��O7�ɜ����;}��2���;8Ҁ�$T5���}C	�e����w�����(��+��/�?��%WV������3�q��78�"_�m�.��+7�F������f���������&	W�o(�H}
�:G�*&g��z���M 2ڭj����i:y�.��F�s��h?;zzԼ:�|���`��gx�}�p��O���K��_�=�#uSys�,�W���3��k˩XE��J2O'���ހ��j*��6�;18��,���5��%����I��%l��z���`F���^}J���q�ƓRm�/_�n�y3	�i�evY]���M�zO0v�*�e��z����3:W�Y���CuI������;�?y�6�{}Z�'�zjl��mS��s	�پ�m�i�Y:��.���?	��[���⠍�{�=���!]`��b)�����~k9�I�gY������$.�e��R��F��ʇ�����'�r����a��q��k�=�/�W63���F���Ls�]�������1n���O�]���7jG�k�K��;�K�Y$��LZ�om�S�;��vd_:
�ĕ���H�I$��г��S.�)���'����0�T#�_gHAȭUJx�)��V
�a�yꆰa�,`�p�P�5�ӧ�X`���z����F��v���}��,0��������#�Lꄂ�N�fu���zЅ�)s����8V���;n<�p��Yq�RF�et��k��U�=�	�^_U��XZˍ��+8��˿C�WH��'���/>�@׻�����z'Mp��!C�MN��������K5
),�-.%Ů⪲d�@�:~R��d�)�?��f'�B<[|w��������]}�m⑐��5zM��z���p����z�F��2}�;�1���$������J'4��+>��c�s1�[yzj�=�֟o%�Ǌ
$�̥Z��������r����Œ7��J�m�xZ�p��)T1qu/�����
	:29���#���a������B�.
s��P�ϐty 7���MY�2���-m��o�ȭ��o�D����$,���~�����`�؏ȡbKd��y��T'���T|�>w�R'E�wp��J,<7�?�]::1����d�%�X*[t���y���ǧ�<��t�d�`gVV5�O7	ou�Un�[��Q�1�.Ua&k��!Ȳ L�Pf���}������ �w�/;t0T<�ǳ�O�0��2�聊���1����I���ʵ/���1hCN�zO��|���r�]&=���8��rt��soJ����I�x�	��
�e�s�RN�,�3�>m��p���VR�9`�ξ21������H7�9.�3�d2L�D��G�����q͚�/zK7��S5X/As{7+�q����&&(K��9Q�w�H����U�i혎�k�q��G��w�O��nU��R4��Z��BEƋgPC������C.s3��X�v���F��w�ڄn�C������[pVk�$WO��'��{���B7?��Ҋ�-?���(/O��V��=`fٝ�I[�0�[Ӟ���`҂kb����kZ�s����"D��N�Z��A�0P��&D�"f�G���Hc���������ުx�'���B՘�ˢ�(lG�;���8o���1�����8��n�D;��ׁ���Yk��?�Aի��]#H���czM4�&�w`
wm4���2ɿ'%���(�J}$�'�OF����(��� ��lc�̓��Ch5%{j���oN*<�:�F�Z�ל����L�b:����	�������s���uy}|���YtJy�>����G��� r	ɉJk8������0�)�N�)�Л ��N:bh߽��x@|�$��Y�9����5�{"�*�&��9���O�7/��|�]�ߖ t]A)�f|f_�ٍX�-8%c��2ܭ�����R�%g�!����/��S����O��6u٪)
G%��(�+���]��:6�M6Q:�Z�q-�R��p��$u�a1 Z�{b�ק=}`c�����0ݒ��R֌m;l{| �6�qw#B7%���)9��댭�����x��?=��<ٙ�U�<QJSH d������Yb�a4���q���s��/�� ���;�&�����8�y���C��xܭ%�^˹l�_<���ѪD=��w��P�J�t�!̩iϹy�U��^� L ���I�C�t���
1��	��'_IF�c0IB�T?�昑�L���ǭ�Х�SE���뇶��{������ ��n=̘���H�{BC���y��ۯ��L�(e�2��t��e�I�*�p���}�� ��2����p�R{�Q5��Ɨʦ��.P�o߸��=BGt�������}Q�b��N��f942hf��*z)�8.6���#�0'��U工�<�l�wo�B��j�h]S��jє�l���5��D*t@����p d���
M"4�J�T,c��0��+P����u�s ����O���VW��.^U�:�"�q�T̕�٭��45}�d��׭��m�'�5'�"�}M���и	-�<���|:=�H�^��"�]x��F�D�����u�zo~�X��peMH���a�wE0��PfX������~��A�����y�A�7?4
��j4�%��U����:�2�*�ƴ�lJ��y|+�Q�0�ڱ�Ɗʍ/�1��l�Y��I�Z��4d�a�$�6�yJ��W6x��(*	���FҐ   v�����t^�.��߇!�	��-.A��j�>�/'>�י�-e1ʠ�WE����'�0]�օXS��6#߆N������)�#å��l��n���,LtGD�.G~�|h���m����h{��}�i8��|!"v��;�������*�p����J�z

"��8��:�yG+�|T��nM��i =f�5�>g7������M��Az�rEx��`	�y��� �|@h��(G�;��'aw����?���;{�@��f�z�f�@�H}.upo�ٯ��i�T�F��e��L�/I$y/�/�����d��3s}k�eEm(�ßv�c��lC���J�,�Ĝ%�J~�A���B�#��Qw�/w���'}������>�{�m��sq��~(;�s�?���r����z3���'�:��+ �Fu�{"�ۊ}�k�)�ڤlZ�8a念��9������Dx{IJ���%�NT������q$�ߔc�k�&��|��"�Q�fj6�7�Ǭ*��Ҟ�De4�O�^�J�"\4�� W.x�n /���B���E�8��h!�����E����Vʐ�tXE$�)��>Re_�u���l��h6j��Q�KtjUG��f�E��%�@�ݠ�#U��)��?�}E���L���a�K&��d���xD*ԑGj'{I�h���F�H_�Q��Q�/��fa�q:�}+�$�[��:� gTU��
s��o�8tT�UM���N���~XL�Z�N3�0��~�A
$s�䁼i}<Y:1ش�d�p�w1O��)j�����i�qc��"*�,0��V�>�9�m#�2����m[��-%�4&=.�!2TC�8�w���9�X�'�菑 [����J����S��Uuu�j��L���f>)�8H�{c����>�yz�
�������;�V�UKA7ZG�|�#cs�z%#|\��R�IBiq�)#A�=�I�.�.�e|$��	�*��
��?J�[�At3�/�� -�@) �!/Z�UQ�!������c�_>G՜&V���&.��o���[N��u��6�;�3<�lb�%]�CI<���5���t�'���/�]�i��vr_S���ZD�l�{�A��q����Y�����j����^ƽ�	�&Z^
�k�s��;����u1�7fA*�|K���~�nS�S��r1��C�[1��Ŷ|�$Vvg��~�tw}��!�,7� ǻT�b�\|��2��|t{��Q���H���m�j���UC) �9�~4oz�+��a��{�3�.T��B,���.���7ϊ��z#�H�@7�ة�����DI⢱���$	�g$v��2�+bH)��U
"#o-�L���fd��ʪ�VK��Vqi.�9�b/$�� ww�C�<{ҝ�~��' ;��V�.��h#֤^�*��q����=�7��!�0�j:zn~݃zuX�m�^|(��xa1>M$?M\=���jC�r�V-W/��Ɩ��ou���c/D��w<�.���o���/���i6�v�9�-:-�
�e^�qP7�������OB<81�j�Q��4���bI�{"��v�?5���czZiy�Qz�?*�v�=+i�e�����OЦ���Ox�5r8��Ƙd�<�W���hI+��T��d��w���4�M�~YJl�z��,Zc�I��x}��o���Y�9�m����wP�͜��Pt�h��]��׋p�V�����&i����<�F1�
�	�j!�jL�@ѨFB�m�s�w�kT~h�������Kh���t2DT���ܤ~�R���Dd���`"_�Cn� (C�D�I�)S��(��Os��ι@�������w��Sc�1�������ŒY���'��A+y+�t%�vz��ͮR��XJ�:˸_��l�f�,B�y�c5��*_���O��G�k��Ѽ�"�]����E�o�:��dg��3+<��� ���ӑ�����WR�,(���M�}��;^�F)a�X�H��'�"D׺/��̱j�nz�}���,�>��N���_�'�(,��s�"u9^��O��mh4[����o�S�1	�*J�b5����Q�w�j~|o�޽��Kg��zYT�dT���6�MO;\�tr[����*Xh1��x$Qȵ�oE��D���].��]��g��w�u���������R��u�e���
zی�9�Q�m>E런pM�#1��c#��s�}�x	��z�����{�:���s��:��L����1p���Oa*��»�.�'ޘ
uVܾ�8���a���"_�=��\�;?k�շg��w� �]*!@����J�as�n[�b����5�V����y�VZ���$BҥŔX;T3n���ԟ�o��S��W�5�g�Z���X�c��+��g�T]��G"�3�|\l�440NNX�q���@S5d�଴4�[���B�����ެ�r1W�uO�����Q_T��_�&Ȋ?a5H�tI�̓�k�@�󰴮"�:]�:�Tr_i�h�>��we���:����L����|h �2�g����3���G�.53�xp?PN�y߽�*�l6|�UنMw�|�}us�d��jh� Z��TV�
E�`���B��s��-��Ƴf;����F��j���k�����j��ƈ4*�oŁ/�:�]0����]��ც��fo�_����'�	���Ͳ�9k��aZ������lL�U;G�@{1���c��O�*0+�s�%�i��^�2Vb4{�i����y�=X�E��`t&��� Bu�F[�V�M����/����D���|TO��z�m��R*9�PI^��w>Ag �Wl���� �$������%[X��`�2�u�f�xU��Ld�������&�,_[����7K>_uV�	�_f]ƚ}�J��|������L7�1B��Bm�D���pQE[۰��|;~�y���Ȼ���}��ka�����t��9������5��ׄ��]� ��ܠJ��@�wf�;βѵ��nOӈO�x�R��Cj�1"|�)$.�Ⱥ/����zݢP�빻�O���)N�*�����U�a�b��3�a���LUs/]�15�i�H�ʸ�DO����j��҈'���G��KWV?LP�e�"{���8G��٫=�#��\��oї��MP;���������o�36Ѻ���������-��;p����ss�<򹸀EF�0 <&S�V�F�-"׺�� u��e����8������(��{�(�xu�G�џ@��)�0;q<<��m�8�o};嘹�&��ZC�Ar%���-�ΐn 9�)}%*�'�4���$�yCP���K$�O�ЅH4�J�	�rO,��#��TPda���vn�O��]���˦���L����gd�x:Bd���Ź��Ě�5ugC�W޲s`s�<(P'��m�GH� �+�5����̤�T�Z1{��n	��Ɗ�Zq�4E<���UO�S�'sf>k7�Y��,_�B{��6ͨ�	O�9�M����.1j��}��\���i�V�N����\zV|����3��pQ�LJ�X��Z\+!5]��ȋN5��-1*/��Z}���=��a{�Te���?���%�_L�U-�D��ej 6�ۼ�f@MaU�"��+�̅�*u4�o|��O�_qo��\�|@�H��]Vdu�ڒG�|���Q�z������ǜ��#,5�֦HA߂IZ�>
���8_QN�c��0���3���hl�(1��n��p3Ǔ��dZom�ž�λ<�͚�R԰�/���`f2���t'���Zъ��L���wg���FB�'W��CW� ~g�)g�� �/s�E[���۵�*I�5��^>�'�ۤ)ҙ����N�q� ��
���<�t�Èp��D�V��hOq��J����C��a��ڛ��]e*S������z���30�L�(�Q�t,���xSkVD�:7��i~���ج��KΉ���fK�N�LOo��Ɠ�b����N����u��"�[B3R�%�qe��殨R�,[I�dO�`+4S|�D/zT����4�0e��	_���`ȧ9W�����,O����!�R��\+�ӓ]d�:��\��r~G�ۖ�:��������u�1W�-�u��J�XK�v늌��F�Y5+��X�Bo�4,f����WXA�Q0[��qz	PY�n����"���/��K3�o�@9�w0��K+�ϗ�k�0!��a��}�(����U������WBẅ怫�G}4�+A4�G����A�O�/�v��<?�	�+ua���@��fȚ�ka�"#QŚ�뷒��2*L��Sb�º�|�GQavt�H�����(:.4�|���D?/v~�\���5�%�]<��;㫛?'�~Iұ��k�(/Jѯt��b���ga�}�l����*x%Ѯcd�,_�O�z'�-��w��x��D�1U/�*s؃���3>��o�q�F�	u>��+F�(:�k,��� 5\Cq����4� �Y���lz�8�g�+�e�30[�ڀ�φ=�Z��*V�o��ó�����~��?�{�HhU'-C���o�4_�܍��\����xŀ ���b���v��d,.��qKv�w�0�o����I�Eϡ��p���8�ޔ7�w�BJ���}���ėEAf-b�f�Ge�����㩒����Uo���#��3���1�.�B*y���w@�>]���y�\Ͱyx%>�:��z<E�=�A@_�WT�%S��b�!@����x�܈a�-�S藈����}�>|��<QK1�뽘+�ɪ�WO� ���pw؟�h��5o�a�D�	P���K�n��q����/�h+-e�'ڄcU��������n�I[������xN�ޖ�B�p9�Hz�J٧'m}w�* h�Y���>�G���ŕQU�j'ךZL>1l�,&F�m��T�t�[�zLA EN�B,x��
����-nwR���䩽���W0����A�SiǠlL�.�@B�؉C�̅�����/OU���P�W	�z�ǵwƴ˜��AW��=�'��a�S#��m����V��~���a�@���ѯ���@�A��S��7���L�VC�sc�䊪�{o�y��]��P<�:��5����j�n�S���n��k3�R�@X����'A�m�k��qfK �ޮ�>�Zu���bc����ex>A�Kc��E��0u�!��,2�Z�%lW�N���n�Aďc}�rY��ׅG���n���R�BQD�ӃW/��C�h4����PK��;࣯���_��R'A����X�����B{��l�E��*&2*�)�)DE�K��%�H��L{?/iH�=GQ��[�b�T���j�{N��G�����Uu9�@�����WutR��+���2R��v�tաs�͖7<܂�; �[������aD�B�x��^����{N�5ʩ��E��ds��ha���Tf1䏜4iU%�}M~����$RS[:�Җ��+~nx�-N�멜QWc��b�-#��O|����~�t&����b�/��>fh	�~b���#P���[H�$c��?m޼H�0�ڲ��a�,���f=X ��\�=x`p�g�N���.3��w�������W<���iWu���zW����Vl��(�u"��e������Ҙt�~�
�̆��6�+�R������ۋ
��'>z|���jaH#�lr�����{��*yA�c��ɧ������V�Ğ~�P�����r�7T��7<�+j*=)EMO���NW8����^Ak!e���B{u��a�m��\1�>���I4P/�pL��n�/�\�(�����Np��8`����H�{@�-�6{K�����=��~�=��X�l<U�wƺ٭b;�X��g���4oliܿ��AN;F�@����:��i<(c��#���hH-׬3&���We��ލ.[O��{>�J�����鈉��A&�8�Ӹ��_��;�k�n�Kͽ���Y�:�o��O�E��Vk���qfe�9��e +F�Z:��U�c�U1�&`�9(�6r8�t�5�]�I\M���tg��~Ʈ@%���'�!�5^��@n്,�u�Wx����t�@Y��DxS���Mm��`P�������������*�H�9��lR��/�=�+�+tK���i���u�Ɲ3p���2�3�C����G�f�c�,-iI��P)�Ç�q'[����:�>a��Q�^;��D&��L�'8�t�=[�/�-lړ22A��5�{�AW:���D.�м�g�g"[�G��u�
��:���/N��>���7I�-mj�X3?�X�.�\�Ǡw wtۛ9Y�e:�ֲާ�"��͵�^��^^��;�d�e�sI��a4I�o��5��7�.`�h���LBY��$�TIV�Flx$X���
"��;[h7�h!�ҫӢ��~1�z<�{7�w�;��6��j)߱���=:6�2v�95�7g���H� E�*���� ~�Z-#���K�>S��N�d�_u�:�D� B��uh����k��X�7�Î���m$	e7�v��b���c���kb9��2�A�����)��~!u��%�}<=C[aTeB��%y�.���(�+����Œ>߆�I��CB�L?c��߲��F�wǖ]���5:\v<ŷ�pI�J�p%g��'��).�~�$#�D�D�w/?V$.-.�����BJ@�ޥ�s
��
�e����ލ-�,Q����H��I����߮3H�y���LB��#he~���������h��Q`���I��;C�z,+� .UA�$�Q?�E�񋇆�J܇��������j&�1�~f�JA�W����r±a���Z�i	t&��e�=���%��N�FW��d�;��#��Í�+�;4a������Z�,Q\�T(4�������[S��J(:� :,����O|B��q�l��76�igXwL�����Zp[������_+�!����O��	M�����"�q�-�o�^Ztf��ϝ�Fsd�2���A~,o���"��r)��^�D�}�{��˜C6כ�-�o�)3��E#��H+F���2j�ѩ����^��Ru�5�6I���Z�>6|Ϛ����/z���7u=����(�r��r�S�|<_Gj�rꚲ��u~�
��/ȉ4��	=��<�M����!Җsq���U+�9��uy[p~R�����e`2��nA��<t���ZYhe���o����v���l�g*�|�
������0�"V��>��*|~��}q}@0�MHό���;+C����M"�V8pߤ�ά�O���T,�l�B�Wo����e�rG{���H=� BDc��8���U�Eׄw{��E+�h�U��3Y�#ƥ� F'���mr��Ke�>��Ɓ�1^�=cⰍ/#'�9B�ܵ'[����m�E�#�	�Oo��0�y��o�T�n���j��-6(��f�}5ܳ2�4XQN�%�bV��+� s���n�@�E��Q�����;<����c��b[;�Li��l��3��O���c?�r-��?����������]o�N�ɭX*"��^��T0�iY�����c}�=^^����_�#G�����Ղ\if���� ��h"L��5,��*j��V~�S�Ԋ����*����)Y̢��,d!����6��/�y����X�0%>eu{}�;g���s�������q�r��x�aiO���"�.�N���Ol_���t�$����,Qc�����q�#��:f���w�R�n�I*	��1��-��+��������K�b�NG���"�|�>}w�1�	�#�g6�W\��U}�S� �[�o�a���E���l�S.p*eұV]Y^b�a�떵{��1l�f�ܲ*)�	M0@ˊ���3k
��0d�z7r�t��v��pT�5^��5�9Ma)�����S�������1eX�p��ݹk�uԨ�NII�(���jS��^�AÂ犚��rf7b�`�i���E�"���ɲ�
�HOYi�����F����"��,��zfEE�� ��=kf��blL<� ,Ql�6Ga��+��ݯ\0��I�\��)|�Xᇏ��YD�9�`��Jj�o�T^�AX� ��=W����W�WB܊죁��#�&1r)t�m����So:��^�-���o�D{Pp�P=7���<��\�%�g�%�d/<�%�`��\�k��2�,>½?Q�?<���B�e���w������@龇]�*���͖���7-�����tdopW��lK���X���蹮�(��Us���p��/��´U+b������U���0)����S�.�׋��.OKY��~��dr��+��z�ݺG�95��d����@�H�͘X�Vz�"9v����.��=�z��S��Uu�2��/l�
���U%Iq�U2�ʎ	��7��;�z���(��ԋ��h��cNǳ�������A��<x�BIJ����8H���c��n���v��=E Ե���\3=U�:�y�z<����]J��p�9��.�:R�iQ�>��fB�e����xJ�����S�V(�$�5��=&B�)Ƶ��kM���,���ŤÁ�Hz�L�q���T�����!q\S�����+Rઋ{Z�)�[k���Pv�ȼ���>W��Ub�`��KT��c��ӳ�O��M���V5^.!2��;@�3���z���F�k���~-H�	B��^nP�!��G��&��j(�I�'�a�I�]��d�U	���04&����L�G\�c�w�<�-T~'N(!W.����s�<�L�**�K`.��\!C��X_�]�ֈ��\�"�r*�\�yf�f�w	}o*�'�&���m�D�F����|��X��D����/Uj����K��s��7ܵ 7�F6-
dl YUl6��z���hqh�.�|�y�(�� ��K�I\۴�6{w<vf�@��n��B�1n�Ё�Uu���	r(#�
y,��V��s+��h�qq7��� d~�S�Jx�C�*�y���N5��S `�����>=�o44\Z������Ű�2��/^��F}�xÿա��5��J��rE�9ˡZ��J����gc���[�@,�a�kV���X��æg]�u#oZ.>�ҹ1������xki��1m���8̝��,�!�߽��E�2�a��FMRO,QЪa2<�{�2�}2��]S��,�����{��~���ȨOy�^J�����*��H |�� ���Y�s�����B�76���  �J�@�8�j*�Տo��M��|�^�㔬�����:@�����紽�)k�sw]Oe$O�y{hy������A����3"�C��ا� ��sY�27>]��g��|E>�l�Q�g����fbԐ�dcg�21,"A���9�m�ԗ�w@��5�c�ź�� ,{sGzb3�$�B�ŧ|E0�Q�
�
�ׯ��wt�*���]��HC����M�N��S��j�Yʥ��p!��2���4XU��Ł�:<&+͜n�˖�+���?㸗��$�"z�t�(���_�?Z_�m:�
ŷ[�%�x�l��_DW� ]5�f>���>sZ�����J֣m�/(�ab��N�^yN��湶�kXϷF�&��]Ъc���Ӿ��@���S�s*���m#��{ǁ-Nd��]�|<`Ώj5��鱜�|ۣG�+�]>�G�+��71��"�FAg��¤<b��Y����]�2�V�,�{X��P��ۏ�VА�y z���_���{e�Tk��5W���0;��9(P�Z������.$��k�;�]4e��G��ؾ�����	*�F}Z�(�\C�%Z�se:����� ��a���3����vA2��`��E�L�����XԖC��j_U� ����>�!,�)��>�O�ּT�Gj<��m૮<J�j���;w�]&������ ,�v�H.Y�R�hI�����j;ܳ%9sP3L�%�[�z�ܠ�]2�����௒������OxķS�}̨�Yc���`+�*�ި�&1����w= ��z�u���eh~�8�N�-j�f���ؽ�5�J�vY�%�6hg��4�'q;�e��Lc���,�-���Y��}q��Ą����z�+F�+َ����Gy�$|WYI�R�H�G�_�9Z#;�y�8�y�W��o�������`fV/ߴͨ��������_�*���M�����o%���s��Ŵ����ڠ��X�������tSL��\��H��jO{ou�.; nRRWQ^2��8�m6��l_azM���]���D�
�*!x۵���8Y�ڂznF-�I�Ğ,K�C쪰9G�̩c~��ݡ񫮍�{?�����Ƃ,��[�n@���f��5��G�>�)���ס2Y�Ӥ�T���;s��~	,����p��T��Wi�ӽ1���uͼ,�y�I7�@����� ����=up�DH���SL��o�I� =&���;��l�^�18��tr7��h���2�dt�D�]:QF��t��O�\N�+B������\{e��9n'����7´X^�3e[j�����V�bs�m��3���H��>�6���C1�j����+�n�`�<ru�E8d
XV��۶md}ia��uZ�����i�7�;��F����NO~��~��x�oc����f�H�:��!�گIO=[S�r#�IN����f��y�m8�N�d��y}7i���j�\Q�YPǏ����:۶�����?�s��"L�S��+�:�i�aOY;YR���P�9�i�=��Y�?�����?l��X����(�oܭ�!���wK��w/�M��H~�k�܃|ى��ꫝ�NX �e)����u���~��Vz�I����$��?����9��ٯ�gc�p}b��	GA�n��^=�}�880���L.P)
�^� ����V�i���[K���ܗ�V�+/�;NlwG��&�vKh=j��8�q�d�3���eͼ��W�nyJ���5Q�zd��a��YI�0���Z'�-[�&���jf�D=`��.��f	j;c�;�A�HJ���{�Q��P�?�,vQ�Rě�!�>#N���u4u��t�����'o��>>$�ܫ���5#"^��J�=������\k�2���M�.��|?R�V����"Y_�*��@��Ӓ������3��G:���H��*��/�D� y�ؽ�ֽF,e�/�-�|�O��]�ۛ7&���f�m"Ǥ��w���tC����l�,�I�>��C�%�T."#=�Md����[�5�uԛ�.�Q��w��� B��zZ��R�{���])�O�ޅ��ٰ	�G{���5UPɪ.?��D65ڭ33��17��lӝ~F����M�a=�n����̎��h���pk.V�="37ߡ�)���0�7� ItH88��q;��0W�a�G*���܃�+�b7D��o��1�/W���Ї�=�)tKd+Xxz���9n��=]�G	>��0�ͼ��y�Py�����Q/꒴{��J>4<W7;�3g֐Hk&�VQG�%^��읚K�i�����2��vb�Q��`z"��api��An@Љ��R�n�OF*�0�.�>l�����]J
!�rZ
����\紐j���\ �.oo^0�2���|����#��q�S+��AM�ƈZL���'�eW�~V�,Y(�.�N{��羂'�I��J�՟J�f�&s��4��H��P�cy�~�iDU�bf2ɍ)���"c�L��r�THڷ&k3���7�B��gVy�^"{�$e�>���$$���65��r}�-P@c&sg��-�+=4q8mn��Je��Ͽ#���tz���/�zZ̞-d|v����'���rޯ���ڡm��l�د��w6c*�p7��)�y�=�3���PY��l���L�B����;�w���)�V�;�ӏ%`���s*R؊ zه��%�f�Hs0e����3q]��tK���ȰI卫��[e�ɑ�
\	�F�x��i4�;��qK
�G�ά����Z 
?#ŧM��℻����餏��e���U�Ȧ�-�*������6���2n�s1b4��L}x��v<2�1�9��>&�i�Bnٮ��DR�h[dD���+���^��-�vѱ��Veׯ��O�#=!z�\ORQ�5�]+�G�=_ll�y?�5mk�B<r	_D��I�L��'y�.�&d��}��)'�N�Ds'&r}GF�;6��tu9�I��PC��T�w�}�Q{����vl(��s���;E�կ8� 6��)�Jq?�_�~L'~7K�	�#�����Q%f����o�s�����L���zRQ��;̋膦U�1�c����|yAl����<;��oY�3r�ʌY5�;@94)�>5N�D�� ��~ukf�w@�������2gt濘d]�w �[�;�3öW��ۥ.�謽��JP�OZ��=�a��3����L�ͱ(Y�*`$��.,�r�1
��l1�]<O*.�{�y�#s��b�avTFF���?�����6T��tV's�a-��՛M��	���[����ڧB��� �B�p̪��6΅�-���I�1������Z�$	��3���@H[�fx*�
��p��`�Q�@���v�2����Z��6��1�1��a�9�"������AM�ҷ��&��eY�_�"�����:J���xD8�p�7譺c���K��.��J�MT�����ɋ�4jx^R��[Ys�=��%��`3;P��H�|M��#[[�a==]�WC�4��@?8�Er3�����U�HXq����șm2�SD�i��֣���Fv���h����,�x4�(���ϖ�O;������� �1��K��|S�hn�'�]��-�|�*ݏ �YweO�U�u��>_�R�"3��-�v���U6Ԫv�4f�_� 7d5v��Kc����Ty���/r1QHcY��z���#�%��<i['9��#�[�*>�ܚ�9+�t=�߻Y{.�r+YSV�i�p3��S���t�Ԋ�?��ʶ6P�!NÕ%���#5�J#AZh�8s�t[׌�����u�Y����B2\�0o��q�76��j��Ab�v�������K�L� 2l+ �dU�U6Aо{	��3�>/�`�K?�W�P��`���1ЍBX���䴄A�V�T��7�AU$ ��l�����*����Rf��������+ʛ;�߃��Cg��'$~����yޝ�\���ސ͸%�� ��H�:�H�W��dn����ut`[7S_�Y�R���K���L�t�"�C�D��d�U���칉�$�&{���K�'�����+�:������5��i!�Q�������s>iW��h����>>Ҿ��5��Ȅ�f~Mq�lk���1����̏)��a���Ԕ��W.�^��(Q�ѡ��7�ӎ�}��DM�y?���(��V�|W(�[߱������O�쵞��sq+ǜ["�2���!�F�r/�
��)]�s��⎀)Ix3"���#��KeK�6j��th	((�P?%���߇݉�frBZ�xMѠ�^��IB3/(�zw�\;0p�� �7K��3�͠�v7-���D���H#�[	
�ht=}$Z�	^^O6؅��6-8ؖwK�n�Ǎ e���\���s{7�����_��7��98�?�n���I������)�T��V��ٹ�Y{�ڋ6_)\�ie�Pi����} _�M	_�A��0t�^��9�ȍ6|*l�Ů����ʕ�1=8d��H����E#�b����v]�|��;Ɖ�b;�1����]��$�)Ux����%��&=���%�y�W�4����V�.�̮�89/�rO��"6�c�˭�CS_��0��VgufGտ����JO�B����i�r�|�gV�;�����5z����P�R�Gº��O�&�4�%�XE��#/O��!7C"+�$K�W2zFM����j� t�sQ���HX���&\���O��o��M��S*������5�q�1�?��zO�=�j�d�ѧU���3�N�U.�ǹ����n8)a�[xD1%_5��@�nY�9�3*���.�9�1�٦SP�Tl�?�9�������s"�3���ҌV���Z�&���c��4��ٲړ�-;�l#O��.�z���ͩ���4wK�U~T>�^�!��g����4Dh���.�~J�v�2y�ȗ�tD\�f	M�%�>x�.��B.�y�`�OfI.	#;v,(���'��䷈5��2s���Ų4�RᏬ�Ng<U+6�T�/�ϟ0��f��<_$�L\m�����1�ӗ�縜+�Z9��E���w�t����8�s���m^֍����+�d^�C߬��k�a����P|�db���=��QY @�?Zt����J�!��02+0���P�^F)5 ��tdX^��>��<Q�)�FX�:CWv�2���e��H��%�]�'� �f$:������~���+�Zj�~x\�rze�s�����Z˽�ޖ~b���.�E9-S�'��l{��X�W�4�lXK	?ĒY���|n�n�e�����}��88�,��~(m?E)��^R�m��U�G�rܹ)�CȾ�5���y�7$u�mʇ�KHT�F^)T��(!H�/�a`�j�e�����P�M0ܻ�Ƃ�������wE�ohf����"�w��6�Cs�
E��^���aB�0d�ei�<~.����1��;jd�H���{���'\���oJ���,O����P�Z5*���;Q��ᒁs�P;#1�I�������D{�T2KBq�ʖi�ߍ�u%]��_�<�2l�E�]����{׽D����gG�
A+�3�GŻ��fs�̏?n���"�K�%�Z)�3�F/v]6�Y��KA�n�\ߺ�a8,.�y��HR~4ѹ>�;�����U�z�h(82�zSb������\�d�8ټ��uC�j.�2����lo�w��w@�lg�cLM&s���\��"_F�p�N���4����؊v�����f?tn�l��.�;n�N�фT�����K^Q�����|8s$��u�5^���OϬ��!�':I�xX &O����O���]�FDǏ�M4�3+�����c�BbۂX�@g�����Jy07�A�i	���G$�\����	��+ݝ2[9�=,����z?9s+H�`�˦��0���
2�N�lF��SM"}�=Ū��3Ucᐑ��}s.��y�n@�A/���[�>��O[����gb�@(#��4��B�	܅ ����c�B����7��rz
��<ضk2S1$��5lgiٮ�0pkxF��(��<N\L��������+��W��d��KV�$�ꪺ;M�k^liˊ[����U��J�+�H999u��2V�]a4��*��&UPj�HD����>CյZGov�gM��SА|��y3��z��ƱȉD���x�5�t����!IѩT1�M<g�u4�BԺ�%$'R���W� N���8�y�Ab�Uh��t��,s�u�!ڦi$r�)�����)��n���k��s�Iqr�Y)\���Ww��U+��Y7H���\���Nss�r?v<#jqm�R��H�j�QT�5!P�<�2~ΕTE��焹����ⓞ	�#Mԗ���O����2N�nC���z>_�A���$r�(D�fK7��v��$�SR'��+��~�?|�Y�3���{�P�=�|�x�����b���?�tS�[�0�UI�xf<�x�؝�`�ecq�S�� ڒν��J����0����#�S7��%4�O��zH)(�֊�����ݞ��5M��r�Y�UK����7�@�?�@f��d "Y�z�(�����0)��Ը�Jĥ23�$Nzˁ�u�/]�����`;��OtU(�q1$�K�vz���Å�sD�B11�9-��dR�����7��\v�%�r��dY�Z��w"ۀ�������Rb��k�6��/?��2C���>�?���R7���сQ�i��h&G�I#8�i,�J�fH�e���E:��9W� �ߣ��C�kLo�G�2y��zO���	�_�I�Z�������IRs��젡 7!/�Mk��Q��%�;u8��v�վ����a�Y�҃\$�B�F�ᗟ%��<#β$#���_�3M8��D��KG�G�Pa������
4g��tj|��I�ZU��i|�����b��ſ*�ؑQzX�O#
��Zn�q����ȒQ-�C��F"���@�����=�LnQ��1Jb�%�����{�Vu�=*P/�+�1��#g����J���^=�'N,p���;zh
���r�(�ʾ�z?�$����P���Rcd�D���D���jr>T�hH�x�c6�KY2�����5D7���ok�7|L�ВiȅV�c^��E��Yc�Eq)��D���ݪh��DZ.H�\���]��ަ$%���'��PQ���B1I+�eS{4q��$���[�a��;�VCt_ "�}O�ާ�{�R�	j����e?y���+�m�g���5�Yi�|i~�΁]Z_�IY]:���? i.�E�_�V��)�	~Tn�`���YD($&�K,a6|~Sg�����5��2���˄��	{�L�`����W����&���r�?x����Z8��)��D����nD<wm���]��*���ӗp%DW�\��x9��4����	��(.^e
�"]F���z��6���g�;@��j��$��D�ٜh��e�V�	M+�j�_\f�8���.��:.��O_i��ٷ6#EU��n�
Z��������&�mװR�tVv���5ͥ� �*��O\f�h����.�#�j�-���W��i���v7�q�l�ۤy��}z2c�o��{tFc�vwS�Ps\�t�N��gn\!Ե{+W_
n?:v2��nڞw�ʹ�D�%�)�#ڇ�Dt���B�V��1����5��$��_aag3Z�m�bkG~�n^$V7��׎!��~NGe[XU�����	E����}a�@��y�!+u�a�X�G�P��Ǉ��[>�gQ�I��-�o7�}܍p]�ݛ]��غ�q;[M�MkD�[�����9c�F�Ǳ�p��AP=L� �z�c��m,��6�9�!.s�& �O1]
��GQp9?���`��?��G��+�\�G��ښ9U%Ta��9Δ��dDkki����L6��B~5Fj$X�a�TV������^�^�0*�1|��_u�E��E�����jlm��Cd,�yi�yJծ��ot�������!�j�DК�c�E|��~m�[�m��+�Qb0�.�E�gĉ'~�d+�bK�SUv?-j��6�C�LP��<{j��oH����zt��'��@1��K	Ӧ[�6������/���K����HVW".� dٕ��.�۵o]H�tq#|�ф�43�' ��,���1b7�_veq&p<�H���5�%�"G'vM��0�v�Va
�C�j���{���L���W-'��f,�Tk����E�ʊ��<s�NzVcs�,��:ò��w�\���I��-L�����8ԹG���H�"t|z�"Ch�^�'y*�m�V�cs[jU�ͭ�<-�U��)�.զ�ZmW�Y�ܸ�IP�:��cJ����~<�
~d�0do:s`>���cU��$�g�AFD�� �/���5=β�[۱S��1��E���NǳыܒAanD9��"P.2/��Q�������a�|i�4\S,���͡��x�m?�P��48l�͌%�H��`���3��.2Az�)?� _I�9|T�����Kh����4��H��F�d3�N �Ce%��W�wv;	k'>�b��Q�u+��x)z �"�<i�idu��D�O�$�2�T^g�yY�|���
��MNh2\�
�R�<����]�lG7%Ŧa<}��̇��K@=��9=�����	�v)��@n_�c�
�y�V	��8��TݒdR����_"�ŕ?����L|�[�Vhxj+'ξu�r^�r{��fe�y�v5�D�zI�.�N�~JJ#X�&�=R�@p0�h\_=Ӟg��.ҝy�/?%��ý��܏{�~(/���h<k剈{���=�	�q啰��%�n1e1�` � EU��u�0 T�c���u-�w^8��f�9������.BMX��%�L�tj���޾z�/�J�*Zv8��%�|UR�@�R�::`��i�������5��)W�-X?�Q�?�BOn�iB��t;s?��Cn�����օ�$N2쌝1�Uܞ�5�tsk���7���dyX��ז6jIx�r����M(qe����8zYd)P{e~�S�ރ��+�'�9p�{V�ʰv`�����+M�x� $��L#���yS_�&f�)}3x=ƂhX����~��#����Ψ���>!�J�`����L�Oۢ�����n�c��>�&�O����UǛ�<��; ���j��;�E�H5��wj�L'�&1?Vw֫ze���m���.������}K�*��_��ߴ��>�m=w�^��
�G�l��?��l����jȲ-�U�{��-1��/󯺯���eڪ�e(���|u1)`W���� �7�=X�Zf�E��k���6����XF�&9W�|*S-�MKF���g P�JA��*+ٌ|Ԧ}`��rT��9U������ ��n����Q����˸E��&Gc,�lW)uM>����5=@�r��*�W�Ƒ�̣�C�$����4�v�7X�׆��B��;k�N�liYv$K�%�`�8���4��(��tm���\ U�
]��+|�|ꜻ>�/���{�]�	�'
-K�;-A��V`�vA�}`�\��$x�J��3Pd4���j��B�ٙ�g�Z�%f��Χ�w�� ГN	�-�Y��;�X���x�=��7�^��~�i��p:�r�y2<�.��m��o�1
��,�\�`yJ�$�с���_:5ASN
�t�y�xO����H��@�2�A\6�{���Gq�� WRRr��C���fR�1�/}|�Y��Qq� [�"�Tt��{(�����������
��۬�m��gF2��W`TD��Y���)C��;��~F�Hn2���\����O��R�m �8U��6{�ki��[���X#�j >!����u�_�>��-э�)�1)}��[R���WG�CWxG^�2�6(Ɛ�3��!����Pn��e�9��8�r�^�a��K��s"1�V';O���/-wV�������pY}�o~�s��ɟ�Fmφmba�i3ی����X >�DT�Coxa��g��!)�#2u��8�i��"n��!:�R�yEu�����W6oQ�-ul��/��v���ճ Z��Z��gc�S������
���y�,mH܎X^u1�g��V��'�B'%��t�1̔ �ѯ� ���@�v�@����"�Ω��Y=.����������ܗ�3%��k����(��rW(��M���8�D��|$�����{��W8[�S�5_��-vLU9<d֪r3 ��aBP���%e1!�n�BrF��J\�Ǔ�$�J1��`):�P	��][s�!��I� "&��k�Rg�u��@�G�C7�	$�=�K�4�,��Y^��; ���P�ϛ��A�m̏��S�f��V�J1��Z"Pt�i�&'�z{J����T5���yIN!K�"�4���-8� �\�8y8���d�ͭR�m_q�I0��>I��T��d��ś� }��[פ��B�h<�[S8ZT����t+;K�V#Φ����љ��_��=�e�}�wj�+�0?��PY	P*n���pAh�dMt|x$44�>F*E��waY�rKx�_��,�g~��&^-g;�}��t���la��nN��4R_��	������+�F+��]Ǣ͏���e|-)C�pu}K�����c��8��P�s��lg������A-["�`hVq�����i��m|X�����)xZ�'��q��c��ф�%����0�S����W����ۛaB* l���w[��Q�(M?��w(�����:+����e-#e������Rz�;��BJ	�%:��1U�Kp�	І+.]K���RCi5q�M���=W����!�^޵�:¢g�9�?���yxy���i��	�<�/�)��I�8��)~���y�}�,��-7�B�}�m��b���w����q����$��]�v$�{�-�����_	�:��=��r�.K^��߯�6�xW���1�G.�տ��C�c�Z�t0����_�E����q��D���vq}�EF��Z�ab�͐�\�3&}򯙡��5:��| �h �XQǨ��?�֐b* ��pY�*���a�]2�+�`�&�M��cx���6��v}tY/�yN3�
����L��; ,]&�$*�������|��<q�i�1�����@�g3�����ü�lY�z�+�`q�5��S� �	���Ab�-���9a�Y}�����L��9�X�FU�m/cs���ЉW�� ���B��,g����X���Ez��Ɵ/ُ:��N�.�ZJ���>-��:�W�lP�^[xM���p\̪N����&��`�I��>Z|<g=��j��Z�#����ƇSP�㢧ː���7|]g�yl��(����"P
/o�)a����W	b'ӗ�>�<u|�6=�X|h��r�p�b��t��x�V-pm=��Q���q��RwQ��dHR�Ԅ�hm�c��T�аB"�j�6��"���S��j�Ŭ��+Q^�`�ѐ.R����$#;�_TAu~3@oa�^?�j��GK�AGW���J'QѢ]�Ӛ����_��K������&b�����ge�:Ft��xm���X���`u1��#��D�EP�����zh��34
{U�h��<�W��`��M����}%]L�+�ʽ��"ğܭ/�y'|��tX9ݽ⚨��3��?-���#5��B���$��Z����D�A��b@ua�R��-�~%�yg���j��'f@�Ka{s��a{�}�
�����is�Ej���S�v��ڋ#d�=���A!z�d��v� �Y~p���g�R@��ФE#�7�Uf�2V񾩜�Ŧkmwt?t�15d�/��w�"��L�<o2��t�;V���͋%�w@6d����ӾjJ͆f�p�pX��ed>}�%�\`�Q�Wd�Aɒ��}���1��u�kz75+E��2�=w+7�?�zc��\p^4:������<�����'k�����]������f	K9b��ձ0w'9�O��>�͟�s,M,����|GlE=y�`��n�R�I�M1�~�蕌����x�v��P:A�l��7���%�����;v+�ij]\*b�!A�irw|��U����_�1��4����?�	����5\YV���o���IV�ߦq���5��i�M�6���Ž
�f���IY� nIo�%�$��hQ �����O�GO~@ӱ�N~�P���Ԥ��΍G�h��S��v	�&�M�a��0�C�E��.�W��v'h3��Q�C�W�&���D��D��kΣЈ4<-�R������z���Ɇ�"��_�Tz<������Ô��ǡ�}�"9W���E���ƍ*qL�A0�:���kF6��M@21�<�Ұ@UO}�q�ڲ����9��9w/Y ���Jx|5�޵�.l��_���D�_����>vw0�4���\S����Ҙ���<ǈ\��Y�qۛ��zo�8*&��T�C渱5��#Ay�Q��`�̵��k���3�Gq��
�Ū�T����z?q���>����4�q�F(c�����u�~4��4N��&�d���V�?�����+�o� H�wѣG���[�w��;AX�*uu��몫��A�UO~oοp��y1s����}��%��)h3���j�V����e�V[s��%���e�����4NZ�ɟ�2���)5Ul$x�\���$u;����k�G�Xs�j����B�Ϯ	��st�}��M?=Vb��߄�LÏ�I�wu��CF�s�1���eڱg�o�A��i�D�Υ�k�����d�9l��&�k%)-i�)��l&�s�-��VZ���������5d��LqDթ���	�r1�R`a6��{�w�����NO��ƹ��w�w��l���9|�W�J���r'W�� �'y�?[�����n�wii5I$��m�Ǻ�� ��{�1���՜pO� �Gi�͢z,�� ��fVua��Z6��]ίI�K�Li��XZ�'���7=�h�S�ԡ��T&������9���u	�^��a��>g�%a�����+��x^�Ņ����>�T��5��
�'�J��M�n�J�;��%/>]���;�!/^�j ;��]ދ3I���ɱօ]����Ƶ¹�����"AВ��!����śX)��r���PL
1����kJ69��*s��0�	I��>P�3]�=��)a�� ���~u����H����-B�Wv �s��[�v/"8im�լdUCV$]iT�]H����R�E3~$��^D�獺�!�j"�H�hB�ˆ�v~��3�Y�B��6�ʜ�N!�\��5'���[����N�-�jX���Yh���������7:�J�a�g�aUU3կXEѽ`���ox�o�N�)+��������w�1E���rY�Va�_������ʆHB-��A�Y��Ʀ�IĄK�z���r�*}O��'[A���"�O�o�pʨ�����������=�8XrV�$2���Y�$��p	�ގ4yʤ��ק�`C��?
̢'�v�_H5PS�������|��?.}���sk0x�۝�r1�F4G�\J�Pߢ
u»���f����4ͅ���&a,I`6���ľ�{�&gy Ŕc2s��nv��f?4�[~����*<->U�T���Q��l�kz}d��:�W��z����g��>Y_9[&��</{;5���wr��>Y*�Qq��oIt%�^������zL�)��)R�G�6yM��s;�\ȉU|rO�ɑ�Zp2����Jޫ	�w;%Ď֒��d�T3��y�QJMM�_[��M���)T��q&��[
�a&�־�C<�����X����w����h�zTtsQ�r�(�4X�(��8z�@?*7�T��������5��5�R^���C���s�o)a��������'������ΩAQ2W�x���k�CPP�#��}���K��C�)�z��<�v��jlo��'k�̰��:.��t�Ւ���p��}]jnq.��� ��Y��T�tP���g�z�&פ���Q���D����7�L_�Ec�kwJE?�`AJS�˖�Xu?E�]ua�c���A���v��~��I�$&[2ۑA��:�7z�)��Ԟ(�e˶�v�@F�)eq?����R�*������S��e���0&K����(%E�|�Y_3�,���R�t��;��x|XM�|���a�$�\W7��;��S#�OT�&D@7��:�.�mո;\��#�@/��;r@�^%�����O��N�������P�U��_`{n��\�iV ��ǃ���}0��W���U⡉�N�#>�C�<�7�P���qF�}����xrh�K�C�&���^�2�����h��r�-V���Z[��s����E<�6�5s�ZϨ�O-��
�FÆ�������>��o���5���Pjɱ���z�����U)��z�A�Z2cu��D6^d��^_?tW���B�p�7�ֿ��D�x�=94u?��ٷ����������i:�}ߴ����R��|*UwF���]Зy+)��n��`jeP���E��?G�����(E#�m��A~���kJ�'@Ty�*e ��!�B|H�:�w���&}����' �(Q�BdƘlX��R'�<M���I���~S��Qq���0
"����"�`|4���d���;��|���8��=R�ӷ�G�a6���=��X!i��ha�C�6�q��lU��ˢ��.hޟ���܉��u��GI�F�D{H��2{7�w��]��dN��rg3�{��n��T�����*�op�˼�GH���RM8|ii�k��j*�l�{��D.���s��>����qZ,m�0���X�H}��/����sI0�};֮��9��������9|05qўp�l����E����
�l*��_f�9���?G���������e�=�Iz%h�:����	�����ꜿ�zu�����3g���BV����m0dW��p��X��-:��\|dLI���s���eÚXdFE�%>BȌ�2�o��I�N:+�@����L���TI��m�9�n�!�l��ο�֖��R���Ya)��T4h�w�%[��Q���-+�-�`��Đ@�is��h�C�Q������my��OPNP��	0P�g$���S=��F�L������'��2 ��MTf]�� +����W�&c��M`���ȶK��Xj#K��I=8��0��Q�eaT�.����-�1��o#��8�l��+��Z�ٌ�c_�sI��8Q�5�
�u�ո�ܫQ6��\<T�CڄwN5�G������q1ɋZ���l��E�yyb��>th��U�*0(m�3�Y��S�|���5]�1PU��8���ز"�D��5RfL��P����d������@�aϐo�\����Y�F����C�թPĈy��zH.V:�ƚ��â;��ik��#�H㴫��$/��t�g��o�\�M�aJf#M5����e��R�]��hJ����(< ����A����7�bSx���������G���}Դ0Ѿ��71�9�B���r�2�����?3�b_���B�p�t;f�ſ���|���!�+���hFn(3I�Pg����K�#�R���_#WpS�y^�k�����	U�����SW��Ձ���e�.v'F��r=�D}�=Q�`רaƅ��*��l��5�����S8��ћ�d���BU#58͠׏'�!�Z�7	��2��?��ZϚ��^X��c⛬0pS�~4���(��1�+q�:�{"���x��f(�~?�x �U�J�����w�2⚼\}R-$� ��^�L�Эz�=�b�`����{bF0�,�����(x͸yܷ�y�	
��Ԗ�AK�Uc�X��:�9bl�D��ؚ�g>���؟^;C�Mz"���݅�aZt���&Ug�93�:K,�50�FҲ����������=�}��$����y�п!�e*�[�8ӟ\֣�o}A�r�i�k��+G���~��K�4ߙ��So��>��U�e���m����w+�^��>1J_+�>���BSw�Y�T�m��\�=z�s�R9#]�_��%�sP�PE�wap��L��3{{x��o<s��v�/��e_I�&&.8u2��H��Z�� [��#� /I�#55�9��B�&c�޴ޮ0��g���\���wNw
�I��c�d��K��ó�4S�KT��cr9��u����[�n�u(�U%�5����3�Ķ��Ji�Fv狢�����ȠG�+�w���*ǅ���ω�	:,k�r�����h񔰔%*�2�7wȽ,:��*�O�ïƤv묔T;��V���X�B�'@�"�W�L�Vv�x&��_�ϧ�3��r`G�ƻ9�x�M;x�������Gsv�����k������N�[g�{kܞ h�;!�����B�������?�su��K�P�l]���Mڵ�WL��'6rP(�|��������ZTY�&&��O5�����$C(O&(g=]�0n�<�@8�G�����3�����^"��|���]�;�rw�'��M���Xk}Z2�],����ۈ�(F��~��)��2��rGb�����|`��T4� �w
7/��ϋ�t��y���_:���2C�a�a���)O���٥�f���dJ���ύ�ՠ��ܶ�,y�)t��$N�5q9}κ��������(�`�N�U���ߝt�;*�Z�|���fm:F��~֡Ů���dS�)��7a'u�_m��,���/H~�>p!�:i��mW��5e�J�p����?��|�Z���v��u8��5rȤ�$p';M@���⟘K��*6)4�����*A�V簜�lH�)�ʷ��r��+SF�zU��&E�'�|��O$9x2��:�����z4�F��}��������	@�uJ��n�[Y!'��/�S����5�PnK�cI��y=<�weX]y+D��&�'������c�7s���,�����
�V.{�ɖ�p%¯�ـL������#��O����	�H4$b��V���u��W�����U)�%c�'J�ֿEm�X��eۈ*�6�U��j��P��א4S����a?T�7q ز$h�x��;��!��W�W�Է�-���x
O�喯p�?o�u�g�Ȯ\��1[�0Cm����%�9��6E�
��^����D:oL|�6���+2P��WE�`��~�	��,j�&ǿ�sUe&&��1�I7M�0�Әt^@���	�!��:]q $�-���ۋ'��8��'���������)��I�������$ ͟�0=��`>Ś���S��C_���:��}�����JMuA܀�$�n��N$ۏ�L9��56�����"�Q4�-��+K�@k�w�C��]��h/�nf��W��%��@5�Ո���5�k�/�cXG�n?��ųfӪ��T�	 �7��|���e���3#Z���@U�D�qY]
M�By�����o��+�/��JӺ*L��+h�zE�>�4q\�H�?��Ӱ�H���K���oc�g<O��Kr1C'��vR���TK�@I[+��es��::ڊ��q
��l[�N�N��g����8���~^�	�͡iYx���Z;�
0|��p����oh�?C)��F����wU^.��[��Q6��IY�1ի���w.�{E#��N���Im}��d���|�0��&����� ξP��C���s�������U��M���F�|WL��i�O��H�(�����z�Ð^�3�8%p��*9�1C�5c�̅T��ʟY���ΐ Z��H��Rܥ�&�q6�����A�4L�4\m�DE������$��I�gy��¹��U��%�F��v�1q� |K '7�oX��:�8�*�0�BW����|]R�h�>��[[:^�:[>e9�_3IO��0�.�K�:�(�ǐ���^��?��K�Wj_6��P��~�
 I>���P�f�b�Z��}����FG^;\�fY�_���&���Z�q���}aބo��i�˭
L�A�G4�[�Azf�S�2cS�2���w^��DK���.�X�c�ݭxkJm��v��5!Ò����W�O ��׊!	=?͉�&y��9f�=џ<�o�ȵ�#%7�s_�����Hb��{��=:z�\vz�ަ6Q=�n����(��)y����:ƺ�Ġl]R6���D��.YU�����,5
=-�A ��"�s�f���ܪ��a������}��5)�ɫ&����z�Nc�7e E|�D�9k�0����F��D)S����)NM����&Y{F��x�iDq�^z,�se�M<f��]ރ�HS�2�T����[G��@�Pj�]���3�����PR�������b����T*:{~���&�����C��ބ.����+�\�������l4��6�!h2C���	��(�F~؎�6��\m����ۀqn�5������~�KW4u�|��hQL2gϦ�������}~���6���x��!�4}_7�j�(Hf�c)���/�"A�
U6�q��R��HH�I�ǥf�2��3:l����w��fq��$̥����(��$�e0���r�D{�ׯ��l�~v�} ��𛊓]�@N����� porGb��������.D���2
�S��z�ɡ��|���f�Q�P�*K�料"�hƂ���N=N^^_���-�P�ca_�i"��=��BY�8+ ɡ2���t���
\E��B1ըYI�-r�{/B��.�� �*Iސ}��Kڄ,t�G|�������YAs�e%�g���zmL�.�F�Ȁq=���F�r�0�4&�G˨Sj���$�61!�[�=8�UkF�"�]�� �ϫ�NZ�I���wlȌmd~w���ca���e�^G^�iD"/�� a��c���}h6�7��E�fi��������5<-�Q!��a��/�Jt-�n��"5�W�'�������.(�^$�s�,�'He(߅�\��������l?:���؝�k��\D�=�@��N�n�Q������'���Ľ����l?cF��@��n<�Kg�W0�q�k��@!M*���W[���l���ɧ�݉�z���:S.0N�~^�V�K��9���-E��Ƀ�S1_�L�Ŕ�9kx��m#��c�{�-����V�1̎cɟ^o+p���q�p^��;��Q0{������ �uP�� ����=��������)���_�K�M��׳"��vTB�3_I�ٟ�`����j~bs���������:��9�Y{<�y��B�eU�D+�;�'���.B/Q&6-B)��7*��\۟~�7T�P��Lj�Έ�a��V�y�M������"X��9��(B>�)�F��B_�pd�����wU��~���i��@; 2�SE�F�EQ��q��s]�Ϳ�ﾽ���xg �j'pTL-�)mNGAz*� 	ʯ�_(��%�u�I|R����v����uw�O�9`��̺ǜ�@�>��[3��s�knDd(!�9t����Y�*ۘO������`��k��P������uu;�͠��d����A5sL����_��-;]1kn14�n^4�#Yx���_�d���J�����_M������~�S�H�3�o0՝��� i:��~�,�5ͱ.��*�'�żٖ;�e]]M�?�������..�ա^{ll�o��tO>.X~������{ǘ��M=���d�[�<�j�Nad����֖'���$��AA����a��=�ߴs���N+T'���]���qW�ʥﺉ� �ZA���i��ո-�}W��I��Ok$���z&��1�Cp�}�P���/�߾��o�rG[:;j��YI_</�I���|L�D��V����k��e�>_����x��r=��y/�l#��ZF��%�.2��{��������2/UM*�B9�u�0Ӯa��s�������S[:x^$���n�Wf|d3:_�{������x|��Ҳ��^ ��h�����g�MX�hK�V�����Z��miy<�������� Yn3ht�Z�f4����G�*ɍ��w�saJ�D��� ��-K�����Iǀy��Uy���2�D*��nj\+�N���@v�����]5�)�n�IN���C�;���e;N��G��I��.}�V�:MF�N�w>�HG��N�Uf�ЩBmrI���R�"{�1-���5�d��8��g�`B;ѿn R��i*D�����	��L������W�?6�
5-�c�F��6���ǘ##�k��A)�iUU٬֥�����"�C/���x���ޅwe���<�g��^Ԋ*������AO�m8yB����W썻�����U��C�u�\��k�.F��M�6r�V+��j񖜟����ً�&F/WYH�3;d�H����x6�n8���Q,�H xZ�r��b��o�0H�p��h���!���M� ��nuM��ky��@?Q�h���� ���u�U�RG�&F �r��ǉ���>���HN�� :����͔�Y˝�DO�0��Ǎ�n+j�V�=9�Sy<�*�,̿Z#r_0n��ϯn
<�N�=)����P˫1�-󵞾(
��`V������V�uN ��e�liX�͟YT[S�m��Cr�,az)7Gx���ᡫ�q��\S��W�Z:*B��^T��&%���' �r9�wGk�� ����i$��y3��ı�!�ġ9�k�b�iD����M�>H��I�{*<
�o9��}�g�k)9RT�r�	�ܯp�8���>W�x���M���d%���ȫ�/F�+q2�C�����d;e�	��Ys�����'��O�ܗ��e�ϐװ� �1���=TS��FUz7�Y����1���'�0E�&���������AFh�޴�KGs�/ �"�h�F����
�2���*}��$���N����P�|P��,Þ'Q'�'���*a[��v�t6v66[�j�wJ��얗&+�c_�kH�ZҰ���H_\W��M�X��ߥ���p��{���b��93������Ů�6��!~�e��RA�2����=�X��vc5x����M}	A�oVE1�'mXW󙊍]�3y��FŦ�E���UA��@I�גvLl���ҙ�������=�-��ލv�c)���L���:g}� �3�,�v��X/5io�p����:��to���Ķ\�ʰ�k��:�HfF�īʌ|�N%$�N9�%�q�:b0�
5\��G�ȹѐ�v�yTt����˹��
���洔D3T ��s"]��%���YW�wIanǷ��c
a|M::������qc�
�b�Yl'��!��s� ��"���j[��)����鼒�&�����"���3�����K�c��B����S,;�>��b��ݦ:~�b~�0Yא��iϝ
�L(�q�R����#��Џ���BM�;���x�th޲;'gtuUqP���)�-�ۚ��pHn�^0��&4��f�@��x���j�+<Y�����F�g���������$��qյȾ���Q���lO'��Bj1GAݿ,����'7���hz��&�.���v����0�Z<M�,�"�`�W(�7�2�w`#��99R@�<wJ��b�p��I?� ܇�we�Z��$�f��ˑs}�����U��(�������q緐+�6�v!(��i��Yw�����|�aS�T^���7�����I��<���ŘR�6SZ^g	$/V��,��`/M����4��;>>j��΃]&C� �t�\~����� �`n̉�����3����<Y�ې���^�=j��"T�xʠ��gR�mɄ���#Z�g�9����3�}!�����˟����e_�����&�K�y�V���,���Y޼��l���\��c�[����v�ݿ=�^=�@$,>xb߭wV^ﰀ1`��"+1ۓs�7���M_��4c2[c
O��k����o��X�-b�>Pt:�ꂉ.оt�Uo��n�i�����̳ ��V������ߥO�����|��+,ƛ�߸�?��y��;67�د>���3Ka������ĸ��_Y��m�W��z�k�ȋ���Z����hǪY���J%�5s6S�#܌~l)	�u�Y�|<~.���sC�
r�B಻d(曵�dĺ��~O{�,C��-/��C|�3#ޫ�Шk��B�M���p���_d��ӱ���P��kO�hX}�އ��Mʒ-����T��~{VJ��W@�����5�����GF��ȍk�s�"m�umm��+hI)-�<O�ZO޼�!�!�<��Hu2:����5Ow����+�G�E~���h\��:p�8˫ӗ�\�����{��!4�<����UQ�L��_�ʞ�[�̶�x���~���<��<�5<*� ��Đ���� j�UF)��l�D�k'V
�"j�>�Nc�E+��l��	�Rs�a_��e����i�͘��LB��n/����'�^��G�}>F���=� @���Y4q���7�e2P����.v��Q����th.G.RƬd�9�MM��Q!�>n������~�a����j�65\�Ip%�|?�5�+�EB��n�[SّhwY�����Ј*R &{f�,�rB�����ɺ/�q�ߤ�C�QwAU�a/ݒ.g:QuLM��&к�#�b�(�R;��W��i��z%vg�RR��&���K}]K7��	�@�(�h�ge��T�DK4��n�2�-�˻��qN;�W�� ���wVZ���r�A��6��X�B��X�	�76����xT���7�I���o9��x�y��g;mUT��k��p�y�E��Tb�!}��$����?�X�����ˁ��;��������Ot��ZE��0��>ۜӄ�l�w�u;X���$/��^#��y��F��S"��;=�|Lr�������8y��dG��km�$���4��y��!�
��~�U����m�oi��nw��<v�G̦.������D"�
dG������ټ�N�R���e3U���=nx�����b#IK��O�y�˞ |);3z�[k��Љ}�O���V��#�ri���ڹ�n��W��8^8�(�J��)`,��ʜ���P�ކ���Xެ;�J�Yx���H��|��<V�����ZN���@�U�|�e-�QTgv
�1�\�;�sm�o�U;İ6��&����0=�qp��=���b���깣���o3�DYm�3v�W�AS}y4�rq[F��:���I�p��w?G+h2	�0�m�е,?�Q��C<�-��-Tگ�t�����w�d'K�aA��Çbc�PQ������Lt�S_	��d�S��'��/#g�L,/(O��>o|}s�5�h|�Z�B�mMDͣf��7�vtڸ����3����Y� h��c�ɻ#+~]�ɸ��~�9�L�$����ñ�d�o6�`�Z�3-�����N���^�t����S��� f���=b��[gT��\�X�
���X���G�ܝ�bn��i[(�W�(MS�4#t�I�*K�>���:��^�kPW���ynB��Hܯ̤Ϊ�!o�y牽�ҭ�3�S�O�
*�\s���q�(��/�f����	k�\��
���L�=-N0fx��s�HaX|2�χB��×ΎWUϙ�!*��� [�%����6�|ωb�C��n���IC��	��k��݁���� ��&
�-|M�& �r@�c�M���պswk;�����60�B���8�����l9^�W-M��c�����Ѐ�gp�s�'���6D�F�R���5S�5z&V񠊘��U3�$�vc�t&-�S=̸�)�HP�eyt:�j�~v|b���jH ��R��8b#��m��Fg��9�7]j�'�R�C��)d$����cl��#C��H;�L������v(e+�eN��>m���]jQ����FgZ��q�a
2�}{���غ%Zޢ]�jX
6��
)��,>,+ɧ��6����|�d��S�P�v�Ξ�VC;<L�O8eT*xx�]�u�o�|)�����b�M�����p�J֞&��D�"1��ڗ�R� Q��NX�py|v���um�R#8�޿y���xE$�C��Z5h[/ �D"�K�ҋ�׋����7�q�Ơ�K�����{_o H`Vf,��Ǫ��*��zq�)s��a������D�N�W�xL�L��S����J�ߏ���`堅���|o���P�T���}��7��JH�Tޯ�����:'�ˎ�P�>�s�%;8i��F��sK�q�����]u�v�����۸�?�[�������(�����綑��*�����]v[��l 5�I�����"�A_�}���Ӄ8��
A�^Vv�J�����&�.Jy�^����©�ϳ�C��Ư�1�]�3س�qI�۹;ַ�TT�k���ݺ���۬n<&,�
d��c�h�����\c�[�/��� ە�<3�a��á�]�]��[qe�O]��<'5Rs3���}X���-��a�q����Ds��{S���]��<4�3�ws��pl��$<�R��B�\�DW1�;G#�F�!�0�.׊pV��0�/�xUba���[5$�3Ғ��y�|�$��������i��\��Ȣ l�����"����H-W�l�7��ʱ�z�m?�a7�7a���y��6�q�}�Ӳ׿u���t�zP�5bH3i��Q_QJ\�D"�;}i0M�P�<5$����.,0L!�=.�v�R_��#�A�������{p��r"/*��	h	�6o�����N)�,��j�w��BJ���l$`�hR�|�_*�}��
K���{�=_�/�w0%7�.��x��������W�:�.�y���P����!,���E�ET�A����k�π��)�2���:��|�2l)i�x�KzI�:��~�.|b�����Hr/;&�h�'��q�t�yINŞ�=?�^��kp���)��@G%G{���7+e�TR|�HW�S�yq���U�"9�R׮�.�q�-Ֆ<�y�;~����mҫ�Q�\����JW�rY]�L���3��u
���Q�L����F��� ��l���R"�/d��03L#���#�~��Xv^��KԴ �WNV�n�ߙH.�|�}����w�t�����vlc�Dog��:��f�X� J/X�PB	���
�s���=� 5��P�G*:�M��{|M�����y��d����k��Y�x�4�9vp��Z��	��d�v�8��4H�xM�"�����:`jqhj�%^b^z�Y0����F�=��H��!ٞs��7��e'��1N�7@၂�����w�����/���Ӄ�;��:5N�o(˷�,�����Wm9�ܖ�E�vjRl ��N�x�F9�EV;�41*����z�VU"�|/kSvb�k׾�&�<�57�AᲚ�w3:A۴Yfvŕ׸�9h�V!>�0����?���������4p�	��Y�j��l�V-}f"�c�P!V�n�Tq�+�wvC���l�� R�O���L���xH�-Z�c>e#���|(������rݨ�����[I+�Vx �G�6j��>K'��+|c���}5=�z���W�?3�*i5�T�CH6y��p?Qt�Ցx���*���*�-��c%�
��J�J��U}Ϯ$Z�����PR����G�R�%�kߘ�ۛ��g�|�q>��HS�7�;��/�+v�����'��N̅Ъ�@�Cǣ�&4��a|M��735�b$�H���9ç�^�[�Ľ��k}bb#6s�R/��|s�v��&nLUʟ`0��K�}ԥ6i���M��7��ZVB?�4�%_�ƒ.�]'��hy���W�m��
�C���GF�C Wdw�T�0C�͕�v�X}Y��#P�����z!�e�ͺ��`�ԟ�U�%�$��DĔ˱�� ������ɛ<�3���pK䃵a<g���|8��WhHr�	P��Sl�զ�C�Zp��m��v�����:��7a��htr�^w�+J39T3ʠ��$MV@:3-��e����:��}�D�Fd_��1dP�z$҇��<��76�O>���'%�o4�o"LN;�i�ձ�E��Rl��Ჸ�zv{�W �%���=gq%7�L��,S�[�������R�J�Y2�B����$���� ��~Az�a���F��� ��%���r�/ښv%IGe��"�D��������wAW�& ж�a��q*o�>��eM���ܵ�E��:�5Ӷ��v�/�gO �갸�Jd�-+�2kA��8�(/K��6T�. d�NƵO5�Q�|gx��Ⱥ3�R(5Z	�J�y�*5��?GK�uK�r��^g	r�!b`��U�*����f��K�Z�)�<~�U��^$�4�
$�������0tzQ"��yoc]v��&��$��/}�t����_]���-n$���P�*}�7��+�ն:�0jn�
�B�	�;���n�mﾯh��f�W�g��^���f2u@�Z���Z��S�W�2ey��7]��XOt�ke�+�`�' A���@��@�X�h���`��:�x�pm5*�v5�>���2��e�V��z��D��ўx��~�$!�x�;y4Dٔ֯�.,,Y�$�s��N�j*@B
�c���<����`Lۼ��q��5ɩ��R���� �6�d�0�n�����m��7�S�� 5��"\�4���]룶�&t�U:�p����<2pCL���ό��]�H5�Ҙw�8��KS,G�zv.|r���[@�W{+�|��v�1����d�,-����9p*;�I*�t��ŉUq���ꕁ�U�B���[�u�sƥ`��G�����:���TQ���ԟGU%��+Z0S|_i��i���A�VVcF�����O�M��4����9�[d�-�U�˫�)�Q�ڔ:=m2���1�_x�r�>Z	B!Û� ,��E��^��9$0��!�x̛����
~F�1�v�丩��F*0Ln����-!�,�7~�8�� q�L�R������5W~�i>�
��`W�,W*���Ё'"�fN\��U*����t�]��P��5�t�T���3k���7-DLjaKzF��'@q�o��Ι������i�������4TՑgݛd�ӭ�GPVVX���>�~��s�މ%��"��iz�ԗ��K�ȬAc@HK�i��%��fo|W���zgU�R�+ɲ��B�L��R����v)T�l]� ~A��q��Ժ��+�鑻˵�?Ј��~"��t�"��Y��G���g臫�o�G�q��������2m�,�%�3�J@�ϫ��jא����y)�v���̈́�S�'�����V�Ep�����S;ӛB�ۦBGG��\��xO��3Jx-}��n��3ԡ�@<f�&����i�n���kK����	𥇙V�~dyy�/l��	��=!+u�B���*�>D'�j՜s_�G�
�1�.Zљ��4���E4��G8�� �d �k;֡�T1ٕ�X2�P7EO�)�P�C�%�=���^��n�z����2����)	�}`���NR�ː�!+��S��N��1}]y�ܤ3l��b.�������v�	V��v�/l������):d�Op �0�P ���:�1a	��}�_נ7+�+!5���dl�sєu;�P�W3ml�1v`�%�I98�cg�� K�$aSQ���Q#�]0h��=��̋�o��nď[�ٚcI櫽���	�Ơ���)KR+c�`ld�.�F���8ƙN]�.�r��'->��󽡬��u�t%����J*U�o�@����' �2l��.��)<\>.�ۻΦ!c+-�ۜ����2����`#�u3Mi��J=�˷�c��m�=�U�0�r<X�͋ ��l��>z>]���w�B�2!���2U\��	5ࠂ˳c�`vAA�N��PX�g8��fcI�L5��^�^��ܽ�%�<~����7����Ƅ��^	띁��aV��$.ב�]Eyfpu
&&�>����`>s�6�¤�]�ȁ(y���G�`��S�I��~�/�)�K�K��aД$�}}��ÿ7�;;%5���twV&wύ���I���-8�Y�]�g��!8�N|��4���P�4� �yőq,�42��ӣ~�g��$h](�{�w���ԥxZ���f����YR�֥8<_�3.��J71���R�|$�l�E�f1)�{�2|����/ń�� ,m;Z������7��^?���֤�h��.��qJ��Ux�*��]�v��M�F�*4�b�֑�v�i��}���o;���8H�A1WS���z�$��ݵI�ş����a����U�辳��%�d }M|�ģ}�6UR��e�W�%��pɀKt!lzʣB0y_rߝ�uI�F;�oN�|_2��q;K�T��6Ay^��%g��t���^U��=�%dӪCj�|����3��-�G���7�eWgKD���(���
�_!����c��<ޚܽ�'���>��Z6&�ٙG7��:S"L��ˉm��՜]�$]���s���#[D^�Aa77��w������A7�A�J}'�r[��T����]��+l��߹v?��ć���<��A�f$b�����,Elx�}��71Dl�g�A�*+�%|��gt��@T�+>��3�������L���"�R�B�A`�{㥸i���'æ����N�ճV�O&�wWD��_�6 �U��z)P��g��_L_T�V�a�p٧[XW�	(�ʬ�`���i&19T�7�e��������8���!A��n�݂C�wg� �݃���%���6��~�}�?aw_����ܪ{O��"���R�J��ͮb�~J�6��j�Ma��ީOV#_��n{h�p'l�Է�e��[[�+��8-.V<�CA�c4�,�w^�������u�\��]��1�]�����"�nY����쭘{�obh�?|و��L)׉"�(�^���0��4�������-�h�]�Pl�����r|&�.� �m�4M<t�Q��1��N����n���dn.Ap��*����E�ͱY�/�o����&�q��-J÷y`�J��'�Ɍ�n�|pӟ�?�����4�&L�r45qx��
��q���7���G����\�3����i�o�V��D~�B�[��5��$�ޫ�d��$���Q����*�a\.��`���x��9Mi����<�ù8�ں�{�O]�+k4aBYaj����<x��p]�v"se�޾��D��f�d[Z����)���V!1�δӀٓM��U�y:|;%��U�p�=�N'��z�.����>���D��*��$5E���M��"��;�����\ߵ����� \�G�m|��Z}'/��ٽm)g�+1�ȵ��<J4h�tl���I|����ۃ���t��?��c&��u?q��st�S8��� �-.si�ZHY��y#��;��o4t�a�n!@�Eʭ�3� ���P1F�ZD������Q�������:ۖ,J��q�\��Y�� Wx���d���Q�~�e��F&���v�7��(ia^����5e� �Ma'�z\\ei�Ӥ`wi��
d��Y��y�-|�%
��D!S9�ٝ𒢅b�n|9W�JQ�m|�M���k"׎?�ٔY���H���#i���Sź�L�Oԝo1DF^:���O�������M��((�h�~�l�|%���k�G��Z;Ҙe(WK[A�u=��ꠃk�g��P�'�}���攕I���	v{hJ�nN���25<Y8)RQM�~Z~�9?M)}>�c����C�Z.U�Ќ��	Z������	�u|���ɉ�NP�2������~9�rփ�����uɟ�˘���c�4]�͹˛�M$�^Ί`���U�����B�;`,�����"|��j�k����oh=KP	�����~o9��ʧ�%��:���A|�#�hnz 6����G��;�����%ʘlJ�Bt���C9a[�K~R��=�g罘E1�Ҕ�rs)^���$������^h&Z�\�|hjXns��u��8g{��V��i���m�?lgȳ�@�:����γl*sl��د��m�N�T�Eu���ܪ�x'd��-��7)˽,U�BΫQ}fL=����]a��@3O-d��ș���@"�S|#�����U��{ҳ�Ӷ�.,�z�߶e������54�zl����H�����6�bVc1H�/1޼oҞ�̰��ެ���F6�A(����lae-$rI�u+-5;��A�{�����7�����.��y�vnv4@��ැ�˒��j��Q����^�V>|�3��!�R6�����U������\^T�d�G%m�d.RZ��Z�����Dh���9�^���H��D�]����" �xAllFFl���9�ǉ�hf�4Y��8Y�χ���P��	'Aw�+R���2N��*��İ *�U[�X�
���:XP���V������k�E�m檀�ث!)�0��
��/��:;L�D��9Ydt���?zU�X3�c~�^����٭�x�;B*�DZ�
��1Z�:K�i��Rp�k���л����s�;�Ĕ�m�o��^�m4�5���c��v�[��|g�OR�ʩ,ɕϣs|��2�^x�y�n� �DDz�P��C���hο�����-Ig����7�2
AQ�Q�>����[W�g��;.��;@{oF6 �����y��nG�db�:쩤&e���
V:g��S5��!o�1���5BM�i&� ���g�'}��M6˃�mgh��f��޹��I���O�U!��,˃BF��xj_������:���udW����&FM8��L�*��Q����C�e��Z���0���i�ܺP~�?HZԗ��w]}��"�S� �����;Q��s%X�@�Zk�~��~��~O�ՉOe�ҜLV��k�)�/׺�*��ِ�7H�#�~���ʐ2����p�nu�.�~(��d��y7���j[H�-۽�+mX�Z�?*)��Z(�x�@A��BK��B�4M��O)��gs��h�,�T>Q��HO�	����A���b(�{D��B]��l���r���BƑ�����"@�7�qm�E�(�/o}	���ikT�����*�'��FMV(�b�s��V�����S67�i�KA�8'l{�7KR��F�.��=��1Xi,z&w2n�i����٬η��B䥲����{��	�]������B]�w@��<���a�����o_YY����s %HMg�xz8�Ŕ�G�=���?VՀ2�~Nr��?����b�*W��vQ��4��V�����)~���%3�x�'�Ƕ�Ǹ7�8��ل}	z۱_�p�L]m�Ⱥ�AIѩئ�#ML˞��bטRJU�B�EsKp\��8�vm��(bt{X��t8�^�bbk?BOSc�G�����Kpn]A!���Jtz�U�C�ǡ#̝�#J``�F>�W�ۄ�RMՓ��`O�C�Q��웙Jy��������Ɨ2獱����k�Ǩ;�CG1��;��°8�;`�̊~n�5ee�kTî��V��K^�iN�/�K?Q�,�>r��G��Z]�կd� o�qyR�v~�������Oj�l� BZ�z�>�Ț�2�-�.�'W,���h�S�-��n�6qvfp�.�����ߩ-��6o�V'�ʧe�A[����_���cYSll�K?d�˧�ה�R�V�8U�5ž*r���[�Ko_�78��0�[_�&���e���5{3������lΪ�[sZ(n�����K��4�G�����[��#� ��Tc��Ι �ŉ[�8�꣡~��F5��s�ݿђ)��q.�q�����|ċ�n��E�!j��J<�/B���B�L��=���!)̈́`�RӟU�ܵ�y�jH�Om���MDG}o�5�<�<��b����;�h��d���y����!�����d=CJ�$�-JZ�5�J̚3Ec.󙱅$�r���s��1��ؗ�U1?�H5�Y����������]�K��4
k�Jx�%�r�]1H�H�J_����k6�j�;�8"����(�F*����2�����#��NP���J�M���� ���nch���_��-�&�C^�s�bē��7d���ĤD��.dg��Dt�t�oZ��ૐ�P�_6r�5������/Ob��y�Y;C�a�9�ŇG�W=q'��0p�%�e�E�I�"�\�l��K����l�*;2^�"�W��0��u���s����9��W��yA�Q��~�["���1z�J���q�s��!��~AU�������SZ>5�>���V��3.F6�i\�d�>���6a��A*N�3`N�i���� ��#-b�"n�C�#M,�)����u�n��P�m6��`{K:";X�θ:kT*[������4�p�]��vz�)����(�le��	0�rr"R3F��5J�D�3yf3�%�c����yly��ͯ��i���J�.>�፽�y�[���������h{Zi{Q.gǪ���]^Kb�Bϊ�/͵��Shf���e�F������R2�s�{o"<BԜ�9���|F��j ��W3��g�]#�T���%}�����:��{��84^>z:j�(L��-d�D�:Rn����y����n���<������Ro��|����Ê��G6�ܣ3��l��$@&f�����1��ۤ<�^ĺ�,�׈H� ���\���|ϲ�nRaR0\�����
��q%	����sةcq_'L�� Q�ok���;�ʚ� �k�bS`��^Х5t���|��*�b��N$�AD� c~���s.���u�ȫ�Q���-9X��9k��'��xh��p�+[���S��e�l�}����5c<n}*��G��֤�6�0�x(Uť�<�K����TW�dR�����a��
�biQ�'�^>�Gvv�es��;L�����/{�m�CO�b���*�w�ނ�ή����(�$�lI߮)�G��	&�dٚ��6j�+[G`��퐽NX�*Q�V%�[��9�m����'�{�?Q(@�rb��"ɽ ����du?�^�ؒ�X�%�+!�ٌ��r�17{�J�p��	�No��@��c��^�έ���%�7R����8�C¤�Z,�ݥ��z,�h���l�z"�e��-<�-e7t�V�f]�3S*��Wh�1��ʈ1+��{��"T`� ��g��8z��_%#�a����hq�.��Ni�`��$��\�U���L�) ���X�5dU��/v>��x�	y����������޾��o!h%��ϛJ?�1�?2���VWԪ5�yH1�z%�K�J�A3VU�73�01�.���b��X@�W�%��"�'U��_l����o�1�][�'/�,3�~� e�se?�ӡһ��*�\�vE��8^&SWkSS�)��	�1eX8c�N������f=�P�#�b�7�}yl��Ù?<pj�s.�J��T���wG+B���%��4\��~y�UrlY&3q]�s�GNB%�S�burp����d�~���T	 ��d���p�JY���\���>���0��ׂZЊ��H���lU\���޴�+xŶ���xp�K*lܻ�a5��q�N��x���NQ4����:��qkYb�h�h �K�,����r�hS�\�y�dcȁ䂝��jⵂ�9�Bj�����xd����Ʈt�o~2G��Ϣôߦ��h�lRlj���q�T��.nY��i%k;�i����X���f���8��v�(ֹ�6��v�9��X��S����)��PQr���]��K@P�n}�z!i"����{��b(�z'�@t�j$��ο�x�R���t�sl�`O�cǩ���@�-y�<>n�)��׷�L�����T�2Ԉ�S��rcĎ�YFq�jN��8�w�=�\y��Ҍ�#��/l�r��Ԁ�cVZv��]�xa��L�Sm�LMCo��eQ��TdO�~���(L��̆�:PE�셄�;0K\�w5���|�IP�!f侙��7�x������롩�S��UH��2۽���X��W� �������[?SYc�#��L;o�7�cav�_q�^������f�����=j^՗�2r2Ӹ�#��$���3fk<{S��b��O#*�_f���Z��YČ+T�K(YTU]�����`C�*8Ov/_Y�:P$ik��P�R̯�����'�\�W��T**+�	Ef`C�}�Tʋ!����A,�i̾�������q�/��h��,�+#D��J"���DwK��.Ҽv�I��mo����_��vhv���'�;�Fg��2yI�S/��Rg�q�4-�B?U�f/�6����p4�
�XR�UL���V��M4L����.���s1�����3�8%)Y׳�/�� ��9����/��-$�(����v|���r�U݉���:�<#�B'���oΒ$��2:Q�;����S����Er��4���3��y������F��ھ��61ږ�o���'�j��;���YrD�4����hX�<Y�R�j��9�  ~'9���}75�g�L
�Lǵ�_jyo��vj�z�y,��b������̗��u���DYICwK�L��>���;��mF�Y�3vCD5�B!β���e�Ns��\�]6��JlY8�4���8 ��B�aC@�t�xm�r3p�O��Sw�b�j�ܧҞ����^k�gQ�UˊVRW��W�<�\�����wֵ����=����;4��y�߶(�S ���=_(������ͨ����@1�o6WJ%���)��I�D�oſ�_�;,l���g���:�tm)�k�`����e![y��M4/B���M_��"h��ǚ�&�i�i�Y\�j/�G�__?* 3>� 0�S���#F�g��.�_;��9�a햯��\��?@���T�1��>
�h�&e�F�M8g��ކz����|1r~|"k��|X�=�.�=��{.�`��Rf5 ��tN�oU����i����\�&�ãҝ��q�]Vgg��bjk�k���=w)��j��?�����/� ����84�M��c,�M+�pi��Ԅ����6����,��g��|���U9j	5u⟭�sD��z9o{f��ny^��{���@�a�8v;U���Q�u��ǥ�nB5`q]M*�?�����L}�,��߸���V�r�������y,�?#R>��5X���T��n�����q(�7Y���Ch\�&Z<Jn]ז���T����=q� ������:�`(�ҷ8����AӶ���ȇ�r��S�nAFʧ��?&S��-���/�c��SE(���+-�I!^%��HO�1s�v��60Y�U����QE�S�Y9�x���e���C}�?�u%�w?��A *����.��u��Ї�0���Z�ϐT�[n���x��;��%���h��)j�7|x��]�PH~=I�c��ڳy�
�2�8F�TҞލvWb��db���;�;���ܴ�t��I[ܽA�@��f.[��Fl}~н#f71�'&��zA�@ui��������ʍ�CЀ��է�m�c�Bs�a�ѲZ}�T� �!�)�:��C.$)�������1��z��b�A���޳yqf,i�4tS"%89GIrӪP��"�����U�v�Q�o�
�aVԟr����N%<o���؟F����{9�;s��u�AS���߯�fVv �����ԯ��絝�C��H��J�l�aq�!N���5u{VJT����9}�k+�f���7A$���ڑTω{1� ��jʫu>;����׎�I*K}MQ@w����؇��~y���|A�Ĩ/y��%�{�/��J6<����T�3+�*k��~�+jk�ej�؋��1wH_�cH1{�[��;BJOx��J�ף���D\��y���J@������7����U}!���ġ��,�[O���f'g�k_Is�kj:�yrBu����2 �S���F SI;h�d�%1[��Z��k 7�<-vڕ-�� �r`o�
}��>f]]�]o_�x�����)�jh�6�h�ղ���-����@OX-��f���i_8+�d�����QȞ�bϫP��uՓ�Vx�~;�	�M����\A�����v�L�b�H���c�[Y<�ʥ4���|�եߪ3�r�^�g4��C�nv8͚�G�"����t�N(c2N��=�<�sz�`�����0����ٌ1���S��v��o��̙���b]�I�5m��V[�&Olzk��U!|�N^�M-���F�'&C��A�,��d�f�fzӷ(����*n_��������b��'w&�o��*S%7e5-b00�����]^�[<��Te�h�xIV�f������	m��\ٗ�gFm����}�ķ�5Bw�����`�s0��p��K�]j�i�1��͇����0�3��eݛ
G@=5��Ņ����6|�ꑹ��/1yY\��{
��Wx˘�t_"���~����U�!6v��lN�yj���*{yʬ�fU���V��
J�Q��Nm1ܽ�ݽhM�ӎh����=����@Lr�V�-k�N�H�\�j��:t?%15�����J�#�2��y|t�x����oJ��0ЯDLܜO�\�"j�met�߿�f�c��-��B 5�	��Jz����r����V�o���Ǜ��̢xN	&�q���X���n�k5r����Q�}�4�
y+�����VR���R�D��vOla�<���?���{a>t�ʮ#p��b�{�G���(b�΃�ɵ��@�ϕ���(���9bǯٚ���s���je����gm.PAv����́�*H��rr�>�����:Qt����-�V�77f��Ӡc�rO��or9�f�r5������e|��Ǧg���5;�'�9*��E�Rр"<�4���� b�>�Js�mܚ���o{��̿6EU2��9�h|f�v'G�h��\��tE����Dv7�M���׉Q����X/5Qw�n�X�sת�pQ�v=Q�槖&�P�DUڣ��}U��m]���;�+�J�t�jo!yt�93g��ς�'>
����i�m�)b�o�8<kG��;�L*V_7O��5�`��A�5�_e;�q��u��8�֏M��� �7`��*�R;'��+��t�S?�(m*x�X����D jO�0аGQn���'�=oqV^�F���$�9[�F�+����5rx��D��S�.�o>.�U� Q�$�(D��6@�H�?s���;+�ni={e��[Upʭ$�`|�[T}+۲��mK�%��bo*����\��!��M~]��P�B�%I��--3KȆ���T>n2L6
3�����8����л��ǒG�����2sm��U��?�S2�P�1P�j���R�Q�^(���]� �<���K�1��7{����3c��~'������d�.a:&B��{�6�Jҁd�ua����b�O.kx�6y��o?��v΁~g9Y��A��s�;U��U�ay�Y�Ɖ�쥔�5�ff�G�ֹe?%�I��ǩ6����|��i�w@ħr��:�������6�G{���g�o��椃������~�;jf._�gn�طb6��jF��.�T��´��:&��8Az��R-����w@j���N8��ؐGT�%�B�W�v�+�2�����5fV����dKg����]=�$dx�K��ӧ��4�
a�ބt�Së?�Ɍ>����~wԺc�e��˵$Qx������=����8�&�S�{�A��3���Ä+�r�"Qؤ�����=�w� ��F�?ŕ���Hr6?�Q���x�,e�l��H�4~$f�L~j���M�TN�����HG��Uh�;��h�_���4я͢&j{o"�Wa�QK�l��Md3�r���[ۋ���Ayo�_�tM�:�]-D�Bm�ƹ����BT5L��P��	�\&�c��w@���:�/�G۪QbO�m�J��0�)�!�0R�,�c�:�+v�Z���+����9�V�*���t;{퍩.\N�`{Wr]0�lN�2q���g�I��@�+�prh��r	����������� �(�-#�v�ե��t�mQ[$�n�'J���7����(���ϡկ�4��R�0l-<�'U�YV�-�s���5C;م�k��cݕ���D�\NWe���&�0[�k;ݏ�j��S��ۢ
6���D!����ØP���:��aY�;�W�S���f��4����4wGFW�?��.�bOO�-�/��K~x���Z�l��P�1Xr�>`�;����=�ɷ�p`��ukgKe�%�ڱ܎���:Y�Ϙ���E�Y����NU2Ӎ
��r��䢏�q�G꾍\~]ĹX_*���":��a�)��v˵i���xhB���~���/�u��v:��q�aӑu�
��yT�q~�����2��ݦ*�1�9W!�_�|h��W�m)���h��E)�B7��q�W���Q�{3�P!+9޶P+K!��@0��~=<��������@|,��F��z��٫���i��~m��V�<�wu������"��3۞47S����u������Y�D�鞢̨���G�R"�ͳJ\���g�+흔�|k#�i��ӕ>ȋzA���������E�A����w��l�����z���p9��P��\�/l�$��5 �TW�+��ېrY�1�� �A��m�P������J��݆|�`b�F�0$3n��p.��0}d+��ث.��$ܶ
��Plc��2����Ꞣ:�g"�:N`iJ���js^�����j�2�Y��ɭ_<�9Ŗ��3s����M��EI���1��g�XȰ���"�iS[1�7B]BOpC>ep�l2Ň����(����Y��<76î�YL���� 4P�o七K���Nƛ}�����@���8��Տ�m�7X7��J�)ઋ��'\��R�{�Xex�Z:�����奔�V�t��|��!%Z���ز<��Z|�vC���V4��S=������_���66;c����ڄ	-;i��&\��c�{�h�Wm��.��1�d=0=���-�Qs��ĝ�C͒245�3r�~��H�3]�q��!8ib��|��?A�:O�Qi�N��&�^L.Lc���<(�4�!��̷w�� (��l7���I���W

��7T{o�m+���x�/�8
Z&�8
$���x3�l��scL.*�� p%�v��X��r���ě!�%u�21�K
�J�����8���i1���fq�.En��cK�I�؀އN#�|�N<R�/�j�W��[�0ؚHm�6j\��=�\�ʐ���
0�q2�����EP�3\�J͖t���d�T-�-V4	�%��B!�X���F_2�,њ��"��y��fC���/�o_@_c�fI�/�Mu��>�b:9ƞ�󒆄���H�s'�/ϿO�|����BYT�x�M��s|�?do"nx����G�N���P@y��F�G��_�o�y*S�B]2w�L�1R�"�slZ�I�8�g{��E.��7ͥ-�f� �w�'��k�D�� �DM�~��+fS)����d�0.�|閂�NNl�HZ�l|�y?U`�p�W�8KKMIv�YXc�?ä;�5�m#��t������ �oR�������R+h�#��@W�&�/F�����ɡ.���_��i�̚j��4���L3�{����uQ��9��y��*����hL�	����F��5;o�g3E� R����أ,�y5� �7��e��H��K�t���7���2�Ld~��n�|��ȐT�(�|���t����1U��f	�aH�Y͞�Z)[IPF�l�yp�������ϪA�?܋����q�m�"������/���80�%���ӧh�9��P�Ю���V�k������~ZH����c}�	�"�-r��t�d�-I�/7"��2 �������s<�"�s�[~F�+�Zצ�����j�����V�롈{B�1@1���"#^>�ςiM"����R'ް0Dq�vO�(�:|=ׇ�AƜ�*~6�"����.Ö�݇�vπ���}�rO��1��{*��86�!��/U!u^����+v[7u��3pf7�K����5���f;o��"!����lQ�`p�u�/ߠ�=�|��s�ך�"���ffo��Ϣ�2_�=ߪ<��F���y��H�j�E��٢黄H'ȣ� pO��>�w6p��J�T�%�Y�2s�E/��z̖�m�sf����F��0z\LJp�h�YX��T�	���7$F~��{i�*�c*�}y%b&��6z���&�!p�*E�oG�F� _x10h-�d�0��hj�P%)�m��M�Y߇~�/�UYܛ�*6��/`j�"��W�z�C�p��_Qy�-f�x4��Z����hc.	5��Y>�Pc��eQ����a���ƍ9DJh�Ҥ	@0����e�w4��*1&�r	� dBU�������QA/2�A���&g&[\
�ذc��%	vQ j�l����,���g�M��~�������/��|��F�7h'jL�t�=�-��o��π��CK�+I��|�V
��8��۴dg)�g��q�I�hAj�?�4��+��.�N�3�7bO��5��w@kiY��vy��3�lS�=����9U�x̡��_�aN)M�-E�h�V�Q��\��k�u���=��c�̛��be�og��y\��%,�3X������V�+����*M2�(���90�JFAnD�O��s�kK��k��Ë��E#wyo��l�oI��z��A�4���d����_�+����7�˥0��\F$(�J��V�(�G�X��cf^�����ϟ2'�(� Kf�]"�@��f�G�ͦF -��W�ʰ��+�W`�����������"��U��h{Gk������_(��A���J3i�j�3�O�{�Y/��{����aaj]&�;��X��+P���~�C_��� iy�j��w����Ē{��K s�s����`w������ʗ"^�xUJ������㯇��k�~�=�)���^��T����C�s��lf��eUj���7�h��������){��E1J�����3�5�!���Po~��]�'��e�_(5lQ,ىJ��Z�L��(��%� (EX���PZ����C��p�0;��f�و
ܬ�;�h6U)�F*�%��o~���8��dj�mI�]Y*���a���b�db�[p�A��P�zm���T6#���>B����4`�U���|:	f�ND����)>I��2���y���������nE��_���1��{.���㨥l��6��ELN��u�@�r�z����ȗ��Fc{�s�ō���&6c�34r�3������\z�z/�Jt3�Tw�+�f��G��P�k�s$��oU���
���?>�u�qwי�&��5�#Â��HpX �~�(�AM[��S�����ˣ��O����I�;��%#������m�Z�|EM}JԽw�J���e�O��3&����BY�������{)�st��{�Ze�a��J�G
n5�㣏�~6�E���	<��'^��"���;��0��j�s��m��fּ����R�T�ƾ�W�t�Ȏ�N�8�'�<�Y�1{���V�m0��y�����6!6�T�W����4؂�� ����i³���)��vԚ�"h���-��_({9QV��֒H�K廢���Q]������I4��Ҕ��z�m�|�j�[�et0��0�{���U$�$c6r?\)>)��������f��ĉ���u�M�'k���d��R�k���M�x�?�4�B|���h���buBMo�Z�TźA�qWn]��q�-��wK̭��L֓Z��ޥ��a�$�(Ď^/����:�j
%פ����{ȋ��V���V�yFw����:t�)��)�/����#����Kr�wK�����Pq0�^^RG���<�1�p�$��?����bι0��
_L4;	�e�8���P��x�g� P��#�䴍�;@4�+N�kc��1
�9�����"��F/\�23��A�e?�[xEX}�7i�S������ʄ���$�-Y��1�X��p�Q�hC'����m�Q	���0�`�q��ɂ�]UZ��[��+.Nrr8*��:S�K	�[�0��� /��^v8�A��-aD���ѦV���/�AY2�d�њ���W���A���v�����͈Y��CQr��t��2q��T��ɡO��DD�k�kH��6���N~���ɛ1�:���\Fft��p�w�����2{�~݉�������K�
�So����Rݸ���&�˰��a��/;oF����6Wıu�-�"�IN��t������v���r��s�E��E��Ge�*<��>�ڪ1�K�߻���^��aF��FI��ug�w��������k�WK#љ�L�ñ+��K}���9��
���j��j)����'���Ӌ�΢�7����c���_[y/��^<ty��q���GKK�q����w�[Ij��H�����#����*G�XiQt�`�H�)��_���; #� VFꋆd�
�69Hh l�����r=g��վƽ��s��t«���{�4���r���y�� ���G�H�-O:��/���ں���G	�g�t��t'�zq��)���>��L��a�к�ɸl/��*��^F��qS�f����4M,tׇTv�`f�ϋ��q�5q�gLߨ���݂���ǫw�ǳhU�B��N$��J���
?����:��|�2Q�㔂�
V&�cr%���D�Vn�a��Om�W�����J�1/�LD΋��W�����}���*�G��l�! ��^iQ������Pp��'�T�|i"��8v�5�EN���T�� $�r�������[Nϙ�,�_.5FI�"�@VUz�m�r�8c��$:�ik�?�P�>��@��٠	�t/��(�&��l⏹9�:U�?w�ig��l���-(��u/���@D&ܙNYh{����c��uRY�rL[�3��}�����F�v����%�oN�>��2��Y�<�9��|�و߲�i�i��Ruf�+���V[ѷg��	D�i!aD�48�сx�����$^@���~fۼa��V�
u�������qD�Z\SqX&�P?���*��mxȯ5�ԫ>�� �
2�7o����]\+lͬR���O��޵7���1a�B��칃�Ł��lh{	6�C<]m���C�Rڮ�"!E�Z�x�_����f��5���v�M��쵡��f~ǋd,��RJ�D�xnH�d�dGMg�B1o�>�u.5�>�T�p g<s�`���޺~ݎ�u�#�դ�[.�� ��1b�?��	�Tr"[��`_=�S0XOκ.�j�B���j �֋���̦ե�zwŁ;��6J�L��S�j���lF�Za$A�JwY����<e�M��6������'Dn��Rق1U����Rz?̡��Ht9����#�af\`V�t����_� �e�ٛ;��]h}��^��5�?�����X�v�M7/��In����G���kNp�ꛏ���_�IO� �{m���q�i�؋��F���Rh�6�q�P@NjA&�"8��9O������eɢ1X�#Q��$��%P�Qh�Kw�2*�y,���<��r�][������ڑ�r�Ņ*�ìK�}H�9gw�+ ��Vσ���I)�=<%T�(���병�5h�; s���,��xz�k�5cľ!(J�Ң�5���-^���v76�@�=�=���i�#��wgP�h���	�/2~#����`���Sф�w3e�'� �O4�b�ԋ�n���s���7j�����=j���)��ZI}$�6�2)q�jit��;���w7�Y�5�|Λ"�9�h\n�~�;್���q��
��|�%4��q�t������7��X�&U��گaV�:9�dt�,y�X��m�����o"��?~9;ԡ��$4�»�`U�+�>r��g9ٿ��+vR�J;ȴ(�'�t�/z�7RB͘S�����(��=F�x�������k�Y�;��=�mv.�"��4����� $��G{�D�����~���Dca,YK�HL�	����Ni��v�N'����:��� �2.���ms��ڟ�#�/�M;�Z��E�J�k�6��7�,g��N|gLF�x�����|$�Bj�5�uO�_ʒu���8��Z�X4�!�b�6/�*��OH�����N뜗��\Ǆ�Q��.x�OL���0�+2��QPo���cG��U���]g:l͒��� �Sk���	F�~U^�1��Qv��pVj��
Ah�O��	��ݳ�����u�����U˙�{*�b8����͊����6�;����:M;ɱE�u�1%�}3JV�ii8�LA��_J�1mJ�b��9�.�I��g{�4d���`J�G���ϼʎҜ�BJ��{���v��nO��){K�9h�9�4SH���ZL�,���M�/Rn��QNԪ��
�k\�j���՗'@JSF��"�b|�v?K���������LF����aSzu����Z��jk�F��{���+w��1���L�*H	7~��+�l|�$�g�)�<���1p��� �@�%-��	���M�@�+2h�/�&`�X�y�π�����[=��1-�g&�-��.���[=⍝���깗h�}�9:�/��y��?�q\��m5��>�E�ˤ֢�i��L�l󺋩q��a�{����
H���+ԅm���j��_�	C|ۭ��>N�.OW��[B��<��:���`�W���"��M��wa:���鳜wr\���>�W�jb#�i���o�9���(���0�Xā=��l�!� sc�|��d����q���q@~�NNy���55��Я$g��j��7"*��r�Y��� 2y�mاG�K�f�!iS7��ec�7.���ᇀas�b���������P�@'��.��kR�O��i��i�}�>4�4���)���Mː���b������H��Xqw�(Pܝ�R��C�]�k��E��R�Bx�������57�ff?�Y����Ұ�2�h������K��ߢ�ԃb+�S���N?�Ge�T�l�6b2�g��C6��3ƗK���A>���*�;�>��B�w���Nn]46b�� WI��馈[�UA�;�{��ΰ>�5������di{�ع�yp~������iqQ{����OQO����F
��?����!A�]�;b�,g��2r�r7�Eg:�!������@��f`�A�Z�o� d�7���)-^�é{R|>�����-7�rcAyc$�Aߞ#�K9�[�ϝ�o�ks���k�_,��ɩP�ګVE7�t'JA^��_���k�rC���l�zw!乜Z��9?�k�"������(ur��i���Y��Zy�D*#	V�ipq��=�R��Q÷�:]����Y
_���8H4�n�]5�H~�]RK|R�wq~WX�~���J��H%���ev������`~d��]�7�;�~g2J)���!LX��?\�:i��v�"�^�W~�z�p�9�)��-4�1�lj�3���s��hEk2zSJ�c�o���T@�Ps�o@!;�����J�$��`y�m �O�����X��&S����/�w���4��10	a]|Lzt�ky�c�k��`��3C?��Yp$M#\�J���~;���|� �/X��J%��[�/E�_�b���J��h��K��J��9��UU���L�V�|]���D�ޑ�\�ͼtE6�`oʟ,�o�?�I�~[7�'?�8I+�"�)M-3���qu��S?Ƨ��,o�^���o!$�ةF�=�Mf��ӧ<��M���HY�k���5Tq��ԕ�ӛ��UJӱ1t`H3lI�{��4�1����}�	�^30�n���.mx�T/���[�ceX��P�}�.����T9�k����z����5Iw��p�Fb��"އ�|VY�w[��:�6���n�����#?���1�M��?�Lԋ�9Y5�(�'z�a�7>y�M~����E�K�͜V�������p�<s���p,BMV�(�*�����q��鶘S9{vņ�h��x:6�	���^��#�s(��ue+$��ӓ���l���Jf�:��3[Dc����լ�βc�����������Y��p=��mL��^(�2�7�k4G�1�׶��d�I���-�� �d���Q\���So[�'�$k?x��{���;.��'�Z�o�����}�U�!�*��,����C D���zm�h����d*���p,��|�zw�~0}�4��ǔ�z�_`Og��.���>����� v���p��$�2����R4Z�
XR�g�����J"3�h1ISdxb�h}ϸ�C���PHk����RN���N�a���;�����y�:��>�w�oa`4�蝚nu+�^+��[.Gvg���G�$G�;9�3|��?�X:}M��A��z�L@���m��,�.�T��xrZ�������[��������p��
SW����F΀�k��j����ɻ�]q��u��E�����5w;��h��S5Vww\i��B=+�=��\6�������6H/k�y�������B�>m�i"��|��������{_ͻz��%I�>'�h9qtzhIʲ'u{�eg�'��"��z�n��@��{S狀������ͮ�m�����4�l�nMmx�:�͠g!w\��9$+��w)Ms�F*T�w��[Rih�)HeHc O�T�C���zc6`�p� >`��+Lh�z�8o;[ur�"���%�IO@�d	.�HKq��ӮHKx����R��-���'+�Q��������U+�Pv����ZOY;�JR�0���k*o㣰)-U�r ґ<7��v��w��0��O�~{C�6C�ϰſ��$WLM���'L�|q�b'�M�Hߩy�������a,��}���W�_�Q��ڶCZ@����i:�!N������R�f0��������+=�;I�6� E���Y���Ӵ���?�o6���Y��3u!tNâ�Pv׿�o��!���8M]=�`sn��@{%�WJ�%f'2��޸�ߚX���u�C~`t��	UXyy���	=�/ v��^�Ϊ�ߒ�g���q�x�o��L���v��r�-��<�srĲ�ĵ�4����S���%�����8κx�\tC��T�M3h�-1*6s
�'%�}��+5����c��e����E�W����T�����V~����7A�OY���X�� Y����7"��,���^G�MI����ĨJ؏x��I9�E1uvp�meO1��?6���d7,�C%@�h�U8�(�/4��`�ܒ?�Y�	�C�!�|�Tjm�ڹj����ĝ��h����j�*��y�f\?����|�e,�M��ȉ�``�	WcN3G�1XDt,�l$�UM\p�[��x�9���?1� 5�*��=��J�M�1�wUzyrB�"q��E�n`5jSqKU�6�/;��}g��;��l�Z&S*?�9�������B$~���M�N΍Ǆ#�&:���[�"V�cq�{�_O�%E|U�؀��ogJq�C���wF�J���B�KC�����6cZ*t�����#&�k�:���?�Q��2׾(��$9ωlw�,.mX�ju�����(p`%�q�����9ڢr1��D�K����
�Z̕?�\j�pH]�O,����Q�@�x��=�C?�wL����ޟГ����R�>��~�߸�+�OV��f �� ���|H�+�c=����E�T q3i*�_ �E	�<��{�5��,���^ �GFJ�&֜o�q�|^es	����y�d�^��3�	r�SB/�2�;:%Q���P��t�����Z�^�p��`H�z��:A^X諘��*a���7���Pͻ�C��x����1�d-��|���H)t4�����6t����W?�E:6[���y�+���Mv��� �M�`J��n�%�S�խ��\#�Y>���n���H�*a�p���5�P�Ǽ��C�~�_���ĥQ�l��{.�]i^?�X:p��ž��L7��'��5����ީ�=�H��	��9�0\j����Ƕ��O.y4��l,qG��:V�a�j��ft��&�����^��q��-� ~�{]K����������f����A"�+q^m��M�ڳ�E�?��
f)(��?5gϞ��z�E#a�F��X��Mغ�x#�X/b��Y�V�v�5z0Ռ���^ھr�ԋ*��
����;�ie�+�a}A R*��SW�`��9z�!����CF��{3	��gg(\��r�w����f$��P�����Hh.6o�kkn>[Z|۾_�6����sR�8d;��Ϩ�H �r�.au� �V��ѥ{�]w
J�1��?U|Ș٢����ۘ��ޯU��¸��mxR,vԹ�V.W��2�Z;�l�0_/hkMs%�b���ѽ�XN�.�U�sU�;�#d���X�}�ڹ%ͩ��IT�0=��%�L�{��"p���!���7D��<JE"��4k�H8��{5�̮�R365�n �������}� ���&�r���U����lO�`BI�`��6\H/��U�_��F�ӝ��� ^�] �䧖�V��ճi�m-eU�B���Ԃΰ1��oMw3��o�IZh��B���ٝ�:gm�@O�XV2\�GR/3����:��+����?ʠ����h1!��=����l����O\O�h+�A5~�p�����,�V��Y��w����2��Ȟ�Uqzu�l,��r���f�N�E���qpJ���Ԑ��L�o��7��f娹��o-{�X�]��jDa��d� W���y\{�X�q�Rt����uu��7���^�����mz��	5l�?U�pl������%Z�/ ֙[��Dmp��700+��,|u"sbI�,�-@��	4� �:Ԭ����$�G��i5y��G���gp�tkeg��dL�,7�܃9��cN�N������L���4�����Fg����V�[�d3/����2˹i�4\BKR�3{�B��N�.&�����@������o���/�S��;q��~���ۋ%�����Ky�-$�i���'ӗ�%RI|�J|M̠�nPy-Ax�?����0�s\�9U���"�1��$��~�����/��u.�KE�������wyD�󈬨�n&*E���ɻ�J��B���E;����:����"�vϲZ�d����P4a�?2�ڜKjG�l���W�š��'���.`����tt���g��y7w����k9+�*>�ǧ�b������ yX��g�3�k�፽ �إ�yQ�פ/���7�7L�#������µ��f6���ޫO��������q�]CQ���.�?�Zs�ߔ�K���xоar��u��Uk��h����e+���9��ۍ�]7�t� �r}�}t���r�� ��M`CMf�H_�p��'.@��OYFN(�߁gh4��>�e��(����^~yWRc����a ��u�{��bg!�������e�lp�8�h?ݐ��!!����4�|�V�V���O�'xm;�s�WS}O7i̿O�Ӆ5��_���ۓ&�}� $|]�a`�]�4k3Z�v�7R*n)C��o1d�z<�t[�ӝ�a��L2<�y=���|�?�
��ٜ�bV�
�^ٚ�G�Dmg�u̗��Ӑr�j�]K�[�H��%ً�i����qu�Kux(�Ƭ37Hc��/2m7ՙ�X��l?���'�?���`�1ĳg%�(��>�:L?4#������%sR�Đæ�H�����y+���S[�@����捬�5NuY��"Y�٬la�R��3֯�`�i��ŃG���?�:o���,7dԅ��%x�#O��-j�$���b�䊔���0��C�xBﮥ�ҹU�5�ݫ�W��Z���1�r�����8�J���(b�&�a�ʱ
V�"f9���@V��s_�<��&(���PS�E]�y`d���t"�< q��j��T�u�n��K���E�}찬VV�۲�K���>p��,{%&ơjSƞv��O��V��,�/��%��0�eѴmL��O="���Q���K����N�{��*���}5���?+�s�WUk�;/�o%73c9��;��;�ؒ�o��T,H�����0m89ڷ�U�,�� D�'|=���3�<�KB��Ó]d�%�WN�� F������י�7�?�	Q�l�L|�O`i�R^�Oa`�h����{�&�ST���M�=  � ��S\ДZG�H��zț����Ӱz0x�
�䏹��Up^ ���~�ГlW�w�1GєTZ��:�z��5q�!�c����S��f��5���ؖ{l�g��bfA�y��{=���'5��nو5w�T�k�1���K)�|kG�$he�յ2�Cl�lS~#y]��{�!�np$�Ȳ���:/��ߙ3�ྒྷi0#k�PzQQɨ&t�����5�>�69��k*Y5ZlY��<�_���J�4�W�q�Fl�|����~��^yXZ5���H!�q���wVA<*�C��#�XuȟzZM�G����Tv�b�d��>�~�9t�uN�H�oo�J��/R��"����I�"�������ZY�J�j�4���KC�Rȹ}M�3Ǘ������-X�ec��gՙTz�����#��i����[`�����$�;�C�O�mv�kZ? )�6�ʷ&T����j����������d��d��,��3��(.��o�H�.D�F�9��S_�OA4^�ћo�|Jn��^WD�
P�)��~hygj�JAX����������B�2�S�T�D?8
Ϟ�1�����B+�m���w��tyט���K8�ع6	�b2�e�Nҵ�JQ��[�jD�d��h�.w������
�$��AO��R���	�	�Ju��d��W���crK⏣��wq_�����:��;e�T|ż.s<1tETŷ��`#I�T�Sͥk+�;-%��������.�Îx��!_5�)g���>��OZE�M��.a�`�y�
����/�a���r�&��Q^����������xǁ�-K�rt��6���ʱ=̕�5�	�/8�gT����ٜ��%Zi1���RL` ^3Q�����ӄ�����;����>�iO�f�S;�+ͯ��S�%���Ȩq��M��N"nd�O��@����w�m��܂���Eus��ק�{����5c����d�u��3���,�7e�>�F9����s��I�	�}���G����}�m���؜�X�"�a`�Ec�#�8 �<){q����k�nG<O�����n�s9:6:J��{b*�J��%�R��/:��Q�2<�6;R���32u��|��j�쭮$��;J���<��*���D��λ@���@,U��d0"�3D<�6�T���(���#v�P^X]�����@�źƸ�'cC�U�<�}����x�.�J0��Vg���7z�^"� p޹��)y�
2�d.��>����ֶJ�(�$̮`�uI3ޗ���M'�<)�d�@�$.O͊Y�����������"n*lZ7�xGوW*do�v��Nādve@a9��B�[M'?��|� +�#N��3�R�.b�X~�J����*&���ǂ��U���%Z���C�mQI��f����MS�`(�h�s��	w��nf�R{�:$�[���+#s�`�L� �_�8�i.�)@R�� $�������-yp� ���&���H��Q�����HAz�>$7� (P�h�x�HI��)���q�-K�1]��D�1�x%����ı���[���&d�G��M�2������0�fj�5��pv�w��E�� ��rն�+C�N�����u�摫l��8����)6X㾺��b���8�N3|W\�d�Sz Hf�����r��0"
����읝+}�����>��`YcSKKW��w�)�L���吺e��S����_�+g����;,��P	w��m?�����l�w��� s򽪳9����;^�t?��>���hN�����G�� l�n��N�����;�?b���VN��M-�L�@�X��5�5f!�����ϩF%�p,��(:�"ɪL�s_�����'.�
���1j�{�W�Gx�����Z����wy�f��pY=�a���n�zf�-*E�~^�53�P�i�m]��s:;��ŕ�(��'j���5a��ɰ�ǰ��k3qW"k��4�/82�7�>Ȅ��0-�5��E ~ZU�ڔ�R<��0)[B�X�ln�0K��/��R���x�pr�Y�X���?Cꫜ�0�^ |_`�����{�rP@�iN��-�Iw��!%��j�^�U��`}�V��?!���Dy��=����`�.�p{E4G���]�j�	�ԕ|����� \�r����!�.s���~�r�I!��9�	[�tl�tª��WB�!��'w���2I���HQ�0�D$���� �w&+U�Su)�4ײ��߾��U���Y�H����SK�rRvH�X��߃���<{�:�fj!����j���2����چ��[mQYЙ���ɡ{��IH�w��a�
���C����d@�����g��R-���"f�W���u])�C�*0���d� :	������lSN;�~�{�LTsO�����G(�Rp��؏!.�h���̌}�rE�6�1#��N���;Jb0Z���YsTm�!?5w����`gȂߺ~ր�\�},�&�2��0ݙcB߽ANZ8��:������ov�����9��/C[]t��o�F�ό絤m���73'��}���1L�"����O�B��T����8?�Ұ������$M$:����~ƥ`�PQ�Ug�/� ]����z��}�2{h�f��ﮠ���t�Vo:[��%
S�n��+�)�d�2²{��S�zBJL�<S��^��hbԱ)¤�Q:rX�×�՚���?�ZG��/���f� ~��H�=,� ^s��#B�}�J�\�d�$4)/*o�Y[�S���6��eU.^	�����0G��o୙��ex=�j���;�'��&����)��������5�5�}�����x�,����2U�c�J�Ŝ7�"����𕸾�j:���Ͱ?}�p����t�N���8����,���%�Q}��!�<��5+> |�h�Mis���Pw�ʳx���s��?E�KŦ�⹨�V��T���$������a�J�ʠG,���=�Z�G/0yc׮%nn�/�^����)M35f,m}��ڷ\1��� ɽ��97G/j�K��rxrS�B�3���{�IC���i�s���i�C�c���O��.�����8^���	ƃ7'O�B	R?KCxb+���`}�Ē��W���cM�ɱ�B7�N�&�u.׶�R%�Y���lS�y��Ft��9�Ϫ�~����(6_�ؒ,@>6{�� �b*��-��7T����=�����2a<�b�s}8���ή��gBS��?��1�iq��߶���dgkDS��\��˲��5ϨP߉Ơl�b7�����5��W� �/q�R|HF/j���UXE��Kip�->'�U&l1����:�i�+_$@t6�y�,��σ�`�LDi*/�X[N/��j���s������J�L���o�#�I��sJ�������h�����}]�?OВ{�~�u0��ƚ�l��g, ��0������7�r-/��NE^ �G��F�	/Xn�t %���,/@�ͦ���5����u��*r6\in�?h��Q��e,ʜl_�vH7K'��K�h����*�4��.)�,�~�dIŻ�>�FK��8���x��'m݂1!�;���J�C*��t���K쬒e�'�G�q���,���m']��F�[`.6���	���YL��&�2��.�������I�4� �<�J�"���ԦL7*m3fJ|�����ʪYg&9������AR�kjuz��t�?1���%�hb� B&1[��_��ͭSJ���O���c�T.F�{�i�)�u{nn�{��{M�1D]�)r���X2�2A�XN��[��K�K��=%���~I��ݍR>�L����LB��Z����Ξb�"e���U�By�����^ҹjל�cj�i��,h�I*Wt�Z��4p����'���Wy�<�0���\ySWJjTt)퉙h���6r�������q6���vr�$�
������`*��"�	Ww�"ҥ����1^���i!�5���/�XAt&��P�V����$b@�*<<0�ožie���W� �Z��aC��hCz�L)΢`�ǉĮ�_�-���
��}r����i"G��5ŬrZz:��[�,��G�j$;�ڗ��_��������� �XL���Ej�^ ����#;�Zf���u��'�	���UX�}os�w�;�'T�}bc�Dm�k�6�J�-�++5�L���B�I*�q�2Ѓ+;;�������C�x���"���]{uh�8�MZ5�5hX���.2��%%�ҝ�_YK#�	PlO�8O���HZ��֌�����{��FPA;�n�r��e1U��p�̍b`���zz���Q�	����?V5o
&1/j��H���T���&�,I����
F����~ �<�2Y��8g�� �a�5m�w�[F�5��E��+՜[�@J�Oy�c���i;��Z������o�uk^�G�T�*���SS���&|kZS�r������C�MW	*S,���}�	N mLH`�GY�� ��3��*e��81$\�a���%9��rL+2�� F��9IFy�<>I���0kgB�'��#$�yLI*_a>�9�)�l���;z^��A7�@��>��3?����m�KW�����BmH�&�X��6�~&���Q]�����E��X����u��RK��TB��M�J\O���A���Z��Z��F�&g��!���c��еgߐ���Ы�@/.����9���e
�H�IIԟ�s��.Bv� ��٘.�����+=Hg���E�ȆIn�FU��);��]���
� Vh\w����ٓ��UQ���+ab����� �C��[�"¡a����ӏJ	4�/�`D�Wރ^�Cc���Z��Ӓ�Eg+�-��ɝ"��8GR���l�t.�iuY�����!!�g���ʥEl~\q����_��-fV�� S!٤2�WZ;0-n�����B�xx-�k�c�=1��3��]��6��Z�h�>l��t��%��li�ȗ���R��,D������\���R�[�U$��	�U~��w���f�r��U�v"Z��s�5?o}�7��.8���jow&�Ce���n;h��o�c���ԯ�f�vsă���&�; �O�V��sa�������c��W��U�����$����{y�J����l����/׆~�SÃ���q���-SY�O��񚻣��}p� �E2���pŅ�_���샿�22f;qo,�-����5���c$ɱ1ѭC�o�^�SA扁�7�4�6�k`S}�}A4���/��C~�)1~\�Pg��E�iwmh�w\[q��0�Rx{՟�����U�� �y,?�'!��M�I��"p�ޅ*8a��找�	�(�C�g,��+��8Ъ�|���m�+��o�x+~�����W�����ʻ�� �O'�E[F�@����+Ex(�Ƚ���6�A�6_��*0�gh��Ę�mo�<ҥH9��E��2������*��R8"R߿}�ZH�����L	�6H����$!�D�m_�����g_��ݪ���6Z����O����+��'*s����[i��cs �<��Wc�������}.Z���?~���VXL�N� 䖐�%�<����Mtr6\�u�ۣuT{0�U]�l��MR{B����ﰪ ��u�U�K��Xo�Ȼp���<w�ְ���ty'j�i���+l�lq���-�(�eŢD��p�4B��AL�����gBb��ήI�������]��^+�a�GG��o��H�@Ig
�k�>5E#*|9�=p�ܿ�MlV��ʙ�E�8��������H
�5%ԯooo���u��w�PR��B������YSt��|�3��A�D�n�� y���O�d�:q�񯤝���.c3M7��mn�J�kz�'j�El�G�
�[,ڥ��۲<*!��N$q=��`�g��N�<��X�pʟ2�׌/ �r(��m��Quǣ����av�.���f�z�=�%�� �������H���E����C�N�y��wV��i�V7�����(2e��]��O=��Q�����vk����\2*C��m�%����5���\����޳�P����ǋV"��'FI[ш��?�7����Z�{C�N���캞Y�c�j~Č(�n�򻰛
3���`f�X=�ّFS'X�r�4ҏ���RN���L�X�`�ݤ��D�Hax�WV>�m�SU�<US�D_����W�#��`�z����{,L�#dP�]��pE�����-�~�{8��9�S�4�6DH����Ψ.�1+;��-7q�<��X)U!J�N���"Cl�e��z{B��W��8/���}��= �Լϓ����a��JpmY����g\`>��Mm(�j��[墦
��Ew�L�� ����6����Ϊ�-�ѫ��؟|( nx���*��vo�G�ֽųg�е�:C�����_ñ��hO,���)w�6�T��5���Qeه<�p=|*������ڑ-�����qS��NCO�P/�j���<��TX��A+�phx�٪��Fx��	WI����7��*�Z�,�,��@(Ҙ��awgs�A������i�	�$��5H��ՇĀ�d��Q�;��Zb2+~�^Q�[����U~����JW�І��%�D��8�����O��
�a-�]�����t����?� �3����#6y�(�㑆��^��S`���d��'+q��b�JԴ�Pf��ł�E�*���� f��I�&t ��8��?75wi��>�	�|/x�)�z���ކ�s�>�.(�����{֛��+ݛ0i`p���(b��c����0DfO���yl/YZ���}��1�5�a5+F#�T��9<�I�]����:
B�(]^O�k9��VX���	=E+2D��b+��2���_���/�1����R�o�F?�Gse��1ޮT']E�_p8�wV���gh�^v�'�gXZ�ߠ��L7��3B�E����0�0��x=�2����B�n�U�����և��jM�o��4�,<u��cK2ͩV �꺤Հ���^���� ��|]�`BBw��U�G�����}*�D�b��,�TK���i>��G������˛��w&�B���y��f;�����ZJ�sg*�^4�%�;y.ڥ���>��A���\QY���&��o��,ZR�b|�U����C\���2�S�'���LI��_u	�W��hX]�����ȯ�b�`e���5�^U'^���ĭ��3UE�}���oò:���ɞ��7��5��/���5�?����^{��)3�A���pU��v�P��"�L������������o#e�;�+���SJ�6Y_Q}���/c����<�$����*ӭn��u=�KO}^��
F*��с�D������;�����`��"�����7���*�\�é9}P	�-G<l������'���
���}-�;U���Қ�R:ew:_�j���̖4lޙPy?��u�Ҡ�s�Ԙ�=������=�
{:������:�W��ؚH��AO�T�v���5	hZ�3o>�i��N1�7���Xm�#ܗ�%����l��:��	�$t-��Gx�d{&tK)��-�WNL�Ur�c�l�����m:�oa�'	Z��%
�����	�9^K�w��rӌ6��C���@'A_���t�����Y�dE℩M��� ��F�b<*���`[�c�.�"�tsmJK��	�	� "�y^9�����(�L��;!�4#h-���RZ������K�V���4/"-��-OP�S��/��OϟK~�=�J,,_��SI���'P$N>/�R��t��ǅ�\��u�MPsy�Eo_ML2���,H���K`�8_ng�a�a�u�b�_A��a������"�~�	yJ9�u�Ni6B��o���Ʌ���t�e^���S�o��t��W�~~%��I'�(��Y
JV& ������qa����1���D)v	ܮ�f�.��v�}�ju�-�&�!�V�|��
�$OK2��7o���J��N�j��3���%Bj�133쵠�7F1�敍,�S�\m�Fa��:����\����\l�V�e�nG��l������5?�(����9�-ؠ��~�ߵ雺%]�{ײ|��HC#T{�"�ٺ�<Y{�ga�n��okh�+~r�eO���z�!�-�U,�:Æ��1���$�PwOt�f��F0�q�Ր9�u2��8�>�H)���@��-;�8�1�J����y��j�?h�<��P���4����r�uX��D�/�j(�-bX���Jf`/�F�����M�D�
� �.D�f�(�u~J��`o6^#ֻ����(i ����03��p�3W��9�\S�5�J(Kd�h[���g,u��t{�s���DT��Gu�,��x�(x@"�Y�DUj
���5���q���J�.�M�wE+Þ�&fטp�,����&�Oq���|
�k�m�sOP�
��Iwm�٩oIc����'+�u�s��{��>�b���|IJ+V�C�d�W)m�$����dwSϐ:�K��1����H����BlO��;{��o��_�O������8�[�Bޝ��ĩ����S�*b�)��!�6s��G�*F	DP�N�aQ�U{�#�J�b�-��2ZǛd��~�N��>�˷&XBB��]9'���#�a�D�[~2ĳ��������P2��?Ki	L�c?62�dt�p\��L�߂�ϱ��{��Е~�B���v���������z�Lmh��iPU��7��9�b��(��oyn
I��R�%� 0iēu��JB��<)[Y�ER%d�L�.�R����(��t��k_*3ZI��/������ aS�=2����2?�%	�ѦU�E�a��r�/�q�U:�����V�,�f��"a#��|`�vQ'gp���[3-?�VʜZ���_��]��[��!ze�|^�&��������9�l��
�-�J�5�u�aro:GXV�W��S־��?���ྒྷ�}5�j�"kJ�պ�q�E1ԔL�_HW8�a}^p�PQ*�
Ht�q�G����)���Kt��x�㝻5tINLQ��E�l��7D��O�������_E�'$����~��E+�k��v$Cܺ���g������J��2��k���a"����l���:��2�to��ڏ_A>q =����*.,�b�w}�|
�0q�9�+��,~����a4�D���np=�@A��C�6`�!Z��&�>��<`�T�'�]C2��t������TgpM�`u��n	zo�F#7�Y�C��n[Kj�\��~��qY1c��m����k�2��=�n4!n�w*3l�s��,�$TL<5�`��(�Ű�2X�`�!�-66�+����z��mV��t"#�=���~���(;L'���.�����
 ��@d�H�Ȏ�����"!gip�o����G�LT�Ճ}s� �ZN��e�V��Ny(粿m;�w�N�+y$���v�/̚J�k$�L��{nTC�����ݝ.�$(�ܻGP�Z3mk�2���Ϸ0����R�$N�d�+��FY�]�o)[���"ϧ���{�+�w��{�n���&�#�sS�R
A�tb"�&��*�
0�y���З?|\~y��9��-�[� 	�g�S���
�
�{,	���sG��yn?2�/ڢё����i֍d��o]֨����T.����*�{��cC˅�X��9,M�E��Hۄz["��iL8?K��Z�R��_0u&���^��,����m��������ٖ��V
��4�<og��~2�gr�`)���TWꉙ�3�zn�x��Dѕ%�u8��_�Q	>O�w����d2qi���i^I��c��˧�}� �i]�ὤО�������W�pC��V2}O�Dn<E:��mT�|�ڽ��T�Ci�AC�={Q�{V$��沗�i�	 n�{���D�qj�JUH��v,���M�'Z��&h|���6���dm|E[4|(�_]��)�G#�x�%�� !�ȷ.��v<K~����w�9��2��md`�'�|�ܶ�i�uof~���/_��k���a�x��R�z�H��/�ą���uMW'+�,X:t�[x���(`��_�E��g�w��}]QlT��}�τ#�/�X����xyQ������`�T>=�xH��R4�Ӫ>����`�w���lGr��؊�;IM��o�z{Gp8|h��@�؁��LwcevW����6q�r7~՟�SY�I\Ş\ ��L_�?�� ��ި�H}�O�=^���������~� ����:��j��B�Y�&�Xr>�O*��[�x50f�Űkƥ0�veh�d�%�!�+�fE�uQH֚��p�{�qfLA#�9Ҟ�L�WЕ�+�1�|���׼ ���]VI�Tb�uV*�fp.��Ee�(�u��S��<�l�6�\���S�vXF���T\�n��Ct�����D�m�� P$�F7�����{)\�#eSt5m����⨕�i�7�mw�|��x11���T��u���$���jhP��b�:;N���X��/>)-�%�F�oR�������5C3T��K�)(�4j��"�����K��V�ƺ;L/'l�����Ӡ�M������.N�?�<+�膖��e_q�h�)>��s|��oq�z�6���8!�5����!5	J2���n�a7q����sC��إV�_t��P���b桢���MC�*E;O��)�wB���)ewCj&��nXFZ������������*��N�nmIiV�����%�:�3b�U��+�C���+N{���}��mm/ހ�?S�0* -�u�@n]9�4t'�4�3(w+XXѭ���T��.�m��7U��5� ��A�7�Q«ΐ*R��)��+$�7�R��'�����Yu��E�:�x�
����[�xq�����@)��A���N!�����;������u��9טs����ey[qW2Rr�rO���!z�`�y�������Dk��%�+tu�=�7�����%��t��B��z�P$�&CY�]jbք��;���i�c6����t!(6_���}�B-~��
�*�R����Kf�=���f �}!mW��!g��PpA#�v'��R��E��o&mZFO��YBz5z�bD�杺��q�5���l�2�`S�v��ٲҁ^z�^Qw/Zx��y��޵=�X7u"��Z_+�,�C���m��ZN���K@�x��|5��t?�����b��U�m��r��iv��[��|�$���}�&.�db�.���ܮ�ʪ	g�z�I�d�/!
�*y`o�{�@�N<�[;�����ɶ!��Bz�l�ˊ�yF����H�F�Yj�x}}p������ݕf[��"z�B��w��k��Vku�l���Iԟ�H[��)K�5! ��*ݑ|�;���x֖!�GZM�C�$R�6��E]�1�ۛ��}+IX�$G�1�&H0�7��� �IG��\]�D�5�$���OuO����M%TJ���E�?9Z#�S ��L��@�0����Kkf�2������@��PP�����_��O����+o^�%)�@0{dK�&���V�g&#���)��[�l�ס��O.�l�tP��p��AA�B��V`;nT���|�R�:&޼���,��s�}�uk�*n�5�i{&$�$A����b�!§�)Ƕ�1�����Bd�f��2Ta�j�Ɉ⮌R�m�?�'���{�V��l*���3k��+Vh(�����E���;j����EfR���4��;����V�����$�WA�ɗ�л�t���ܔ����t���r�DA0;a�� �-ˣ���%f0�vAB]f�]�;��F�p�rj�W��HT%J��G�$}g2`���d� ١[�".�Q{O$Ű���1���`�!����*�q��\�/Z�ܤ�fG�zkV%�*I�H��胰���oR�ʳ�U�G�[lB;�H.mN��@��H���$h�Y��6���E�K�֜m<	�Gֵb��w>��3"GQr�X#�H���bq/J �Ba��b,�h
�CL��{�C�p��lֶr���ʰ����S�Qj�0�K��J���hd��B�4&�@���RR��2�Ͱ���Ţ��7�{����=��j���'�Nyg�+Y�.�
;���R%�<���|0�R�kv�����h�sd%3����{�i�d@㌼n�\��Ϩڴ�v�������42��W ��������N��д4h�[s�c`Tg��*9]҈8��^,��9u��0��JM�����\�c�l��KOi�;|��$&&��{��̉L>yu���S᫒�9�Ce��ڋ%|p����w9.���U0B��+]������´�xp�y7f��<���$���C���O3�ɸ�\����΄�4��LG�Z����r�̿�|��k-�3�� )q%�3}��K0�A�.Ŋ�rQ��j������~#Jw'�ԩ�y�����3��w��WMh#W�PPf��qil 3P��QG����|T��t��-K����=5dZ�q|Z���\&T�1?��jǉ�-�
�,�����j�T\ST�I��P�}n&:Z�s0�
�6�=@�K���b��t�+BH�ݹ�-��6"��5�6����2��J�!�B��������L�[� �ȯ���ټy��?�OR&� k55`�{r�3DI��t���{��:�W��,���rxv4��l�Z�<�G��1=���<G_U4���P�_���C��
�)�q��Ï�q��T��,�!��Ϭ��/m}5���b���K�	��}^Y=k{Z���p�wo�]]h�%�)�\ր\�xTHE��I*�e���D�r�VZ�-|o�������`H�7^qr�iR��=٬�&dKG��-��^jʴ�F9l�l�R��u�.Ҩ��S��^�q�r��cv^�u<����A�,��2J�[����䘬q�{���RAG�^�x=CA�C-K&i� �4<���XVv����(�2S	�ů�!��E�RRR�3ټ�������1��5|���grAGT6t�b]G����dJ��f���O�f��$��'�]����*y��Y��*�+�PQ�v2�/-_�� ��@���-Ww��h�-�UHT����#.���ȣ��Y���j���l����c��1q�����oz�}o�����'H{绬I�r�"OYB�1�2��j],�5]�n�n���6D��Kj-�uC	�[20��c@�?��H�����{�~;[p��4Qeޛw�8��Y(Q *�)���͢�]l������(e��zR����.��(g�g�?;�.�\������Z��^Jrg̙]��IJ�r�DQ�����!%��G�g�X��%|��JW6)|ޙ����t�N?R:m��4�m_&%�`o+&9���)�)��¤H~rUzܔ!�	��'�e_��s��b5Pc�譛�0~���#{���9���$<!��ȋ��㒄­i��([�#��������)&!�Y�<d�D�5����Ik ���Ц�G��M��H)�;��g��W��ww����RH�C	�2���`6������x:���������]R�����������Z؀7�o�v��Dp��U��V��1hyw磠n{�j��0@ĔŦ/�;��D���dl)���:�.��y�1,MA�3O�C���j47wP:]��%o�<�0���CJu�>v��E�F����.ݐƎ��b%>��MA16-ى�nIn*��n�I��S��>W+�!����.kٖ��@��<!�^��4:��o:D�����������+"���`E�#�5%�TtcQ�c��VHs^Ô�����F[StI�h�����br�x�)�M�0]X���)ì㣓A'|�g���1��!�Л�6�H�#��<��V�$渼`Ƹ����]�-��

���'��9/y�(g�▻�e��#��q�����
C���,�y�Nl/f�����
��ɜ�u9�xN.��n��<������M������RXKK�^����R�+B?��9����-��+`�Ֆ!��������*\�:N�{5�+�����xt�6��04H�֘��a�
Ș�4�R2�8�c쪓�S�inp�~&�H�4�I*�����x8�Y���"�>��C�^$Z�b��B���_���MBTs�@-M��6w�H,���G�hvX�*�ê�Y�@Y��k���H��l߼�ot�?��e�-��[���+��M��iԺ�	�-?߬��s&[��"���e]z��C������p�>�vp�g�v�<��v�.�^.��Y����Y�-e�  ��R�׸>��j�U�N�v�T5��I�_�~�=��nݵ����X�������s�=�8Q�f�G!�QB[,��uLF@žy���쀮R��V<����-�A��N��,^-���vBe.��U��xf�ٱ�"
�o�:���z�\�Vm��td���F2p��kn9t׆ۮBVO��D����ArHޙ�	Q�/õA�*I�Oۡ�=���V@�����YLE����w~��d1q��z���w8�*JX�R2�^�Y)���eMN�q�K2ic8~��M1Kz��QĦǈ?�=�]����Q�VdUf� �XY�sq������[.�6�P�xx2��h��G����\i��hg���0��S�P_]ʾk,O6��-Xb*W�M����}��H��P���+i��n"G��Sq_�/*ı�	K���:�;ee�23�U۩U-:'t���(V\jaقi���C�.�������ZX���8�Z���Hn����G�F��,��~6��MF[�wK�Cļ��x(o���!�	�6�O'��kKʘTF�S���\IS�Xz���!*�jdW������u#{�ӈ�׀8&.cQ3~��G�F�w��L%���eS����۝�'U�WF'#B6�\���>�Lڻ�.�G�6��*2�X���,�N�	���n/�5$h��a:0�g���]M������D�X
��B�~V�W�U���s�U��� C+��*��Vu��{-��\t��ւ�J/o�"�
���Q}�W3�
o��2VO�DB���/������k���7x<�o"p���n����}f6�5��9���զ�W�$�>�K��ZY��ۖT.�Ȁ�R�O��*	�6�\�����*
��H��25N��T���g�Y}�QQ�>�~�X��{��{kbw/hO5�}� �T�;A�i]qXhn�o�9���ݡ-���N�]�#liSD,E�~hz�3Цh;b��3?�xs��Q��O�n�Z
�Ͽ��R��E�N��j�QD��qq��_��p	fPR�wt!�܊�:����K�Ma��'�Y�7A9�
�f%��3��i�B
@�E�����i-�S��R�����֐�����gޡ'%R�\J)DUW�8��a٤�p��Nb�E9olhp���M�L��#P	O�CJ�O�4�߯��I�	*���"��`]x}YH� 5�j�S7����-�œ}�-�u�
��f�����"��%�<�)�ӐJ� �F@�S �-�b���[M�O��	U�Ga��i7������df�m��I���t;����E�h�0� 7�l�S��w�&�L�M�?��&��7��<N�`/��o���i��6���`�-�fY]7W�8����e��X��(QD���fr��-݋��Pԍ��:�����I�/�b�/f������4&��EL��',U�;25ce�ڡ���]��N�Sm5��[	s��&Zj���x��ۊ�d.ML�F��o�����xp��ݣ��4;/9N�qb~l����B�����E���n�x��P����N���g��ޅ�è��d���B��̎�{��l�{���p��3t�?�CL�|�:��Y-dR*$Ř9��9酩&�p=����I]5'�� h�Y�i
I��]���{ {�h���A���s'G����A���j�y�}�w����ú\��cƭ�('*����t���l��ж��	��b��Fk!%9�inU��Տ%v~��ê3��7�o�ߦ��<m�k�e���G^����2��5N`$�䎽�-<G0��q��������8�9���w�ݹOa�3"����6�}�)̺V�?wO���
�s;l���{%*I�m�����F�C�V��KV�X^fQ=��(�N�P���Q=6�+�JZ�կҩ��WE���4N�%��tn4q��C��soztὩ3Z���&���s�����:���4\����
S]������<ΰ��X�ӓ(�%@bw�V�	���oaO����yKօ��gɷ�;���= ������|Snxv�g
��m�Kd�4�yIa��-3g��8������$�=!��@��c������/f� ��=\���p��zA�����V���������V��r�h��O\>X()2O��^#�wp�)�N��������5FM�	M;�M�����<	�Vч��ee�5��4�
o�+����y[
-
R����ljU��=N�kS�پ�k�9�3v{S�Ee���j����	�V�și'!���͑�����$#���S?�u1�墹��f`8:5�W��X69=�/����+�N��q���5�:@��'T����S`��pRi7B8�CO�"�'	�lÍ9"��]f_�� �n)�X�E��
���^�@�L�#�갳�6����v[��͸��8�D6A{:ᵈ�V������U����8,|�u�~�8
m�DJ�lsc�k__���p�4M�
��7���������ky�Z��2�>�1ٖi��͉��am>]���6��&&�*��{�c,�$,����<��O�ř�o�N��_Y���xe���}����x���ViPS��,<la$H�^£qH��ֲ*h�tʎ��'�~���i�	�\��L��PѠ��c��1at��0K�[?�|Pq�p:�g���|��8�)�3�#���w���eeOJ�=��k-�\����Cd���uh�G�}\��*tk���y	��㯟ȬL��zr�m�T3qqQ������(T���}ŷ��9G,�N��e�/��O�h�?�������IO��#���J��A���&�usM�ϡ<���mn�S$���ؓ��g� ap�K��g3B0�Ǵ�F^H��	oW|��Q��i���
i#o�4ѵ*���M$���Y'��O�C�_.��E}r�j�xHkr}��B��L��Y�����وra\�,������=���l�o����@e`�m_bN$9R u��N��ʩ����ޔ���)�N�s�=~�K�o���.Z�K�;t�u6;�*Y=�7��?�#_tk������6
��Ú[��x���P���Lܵ�s�6&5�3J(+t��
��QUoԲT��B�1;Thȩ��Y��Ќ��ݠI}Va�2nf~�&6sZ��'7��6����[Fb�S�Z	��"�>�H;�`��ݷv6�8�µ8=+Z1��Z�:*«�9�Ű��@��>�[���%~'��xm�^K�� K��L���5g����aS�t�媎��T\�T��(��_�=�_�]1mm����m���NO���2m��>uvfCN� ����E���LW5���o��֕�ݒY����>p�y{?�|&]j��e4�a�E���(��"�������4��9ɿ����x��+l�;sp�b� zX��������X�3�5�e����*m�R��?����ɑ��'����&O@��O8�$��be/�����y��b�����1�������*M�Y{�"��I{~���P���Мrc�B���Ni�W�A-~5�S���?O��ld�� ���U�:�'��Ԗz��V����RD$	!Ӎ$(^�:Uӯ�t�/]�l7p�t.�N�M��u�/J�O+��r9ەp�bWbY�8$ug���Ա�\�����]��W �����Ȳ���	,����g�a����b��SL+9�W ���g~�\�bs�i@�O��'���\��I}�H�6R� �"���;�* �~=�?�s^��g��G�1��昗+���1Vȩ|Z��w.#���l;|�>��5�a˃%�5T�N�����Co��l�vB�n6f�xޠ���w�Z�c���͇�J���o����6]������60Wӟ���d��4����4�*��H�OBG�*b͆��[vz��b(*p���>:~���^����֏p{ӸM�m���!���}�1�\^�?Y�X&���lydZ\^M�Ց��w2�W��ݹ�2	���jpKPE.�j���V�b���?�P�u����e�dp��e.U�[���Y��|�ϧGd����A)�{*g��ƂU������3�/�d.Y���$�Yy݋�kxC2$L�Q� �49H�����ý��a�;��z��E�=r;��=����bO�����s�������3}�R𐼴-�
��j��d�ݺ3�_�?Rv�
)X0�M�+ģ�z��J�����>�:<S���/G��o�2`;�:r$v�/6 ��[��V�=\_��aN�����7q�[���ğ�{K�1�b�g���:�-�2
M	���Bn�o�Y+	}��5�N�q˕d��<B���f^�=<7 ����k��u�Ƶ�[�!��Pu@)�f��$#2d˪� |���i�8'��`f)\�U;p�3�60�����xY�<=2��n��5��|�H����UQ�u�̫��D8%����3;���a1�tȯ�C#
�\#ى�PI�t�J�;y��B�<B�F`��"+��w	%<�Rê��+��bj�6+s����[%\X{�B����_��eʗ_~2&,��@�|d�K��z�:�c\~��Mu�c��<�P]���H�6�J���5�(���"�oM�ݛ���_UL�
���UOo=�c��.]���k�e�>Wy��z�)
����W:����=���Ѫ�
/�H�e�)�N�8ӗ��fTI�} Gd��.�,6���<n�����:fg#�;M݌�&�<C]���'9�������ә���٠����J[g�ŝ?֏�=���R�˲x +��.;��ح5�?a	,d��d��q��;�ok��W�O����
��}"��Ψ&&ъ�v%�LNF����]~3�9u܅r_��_lezzzۿށ��}�<��*>)���i�5�䑇h�Uߥ�!���A����N�Xt�75�'�.I���k��̧���e)�8�3t%��H	i4�nc�[��
H�Fuy~p��+�?���ݪ��󍭺Z*������������En�iTZӸ�N\G�v�]%���%]3��-&�e���5��7�2�ߋ)�B��<�j�x��3��yp���|���~��� Z-�B�R�>|�메��2��}��|b�
�2���ċ�A���e�e�%�v���_�H����H�v^T���_,����nn}Z����-�W�!�?#X��6�g:۞����D򹺆�~��ɫi(J�<��~g�\fa�hj���.�@�ΒM��a��	.�m��j�D��C����`�A�`>1Q���/��p3�;m���䲛Q6��N����r"����lK�owB�c�����~�uArd���zv��uE�`��>���?��1m�m����r��8.	<��ş@<���#���-�Sm�nŗ���uר���
��^��F�ǟ)9З'�Z[���V�3�&��hy���e�k`��I�ڸ��������N��S�:��Ȥ�H����op����n�7��x��,;�J�Yi�yO��ny���I�����ޔK�I�]w}oǭ]@�:�g�H����p9)b�ة���ȴ<D�)�͵�%�[;J3Mݮ^La2�rq����	���+��VSBY�TY����Q5�/6�c�Ū��Hg@C��M?B��>��~0�`�Q����b�r���欫lf�z�����[iҊ
��:�˩4����Kz\̥����32`�H:CX%�%��$rheQݲ3�J�� R��!N���o�KdSsr/n��[��f"a��۸�l�G�cl��Rg� ]�����&���b�1��q�hJ��a�6^��g�C���yu'2&�hx��1�8��AZ&y���6�� ��~�
���v�����-9��;�y�-aG;f7CQ�9[,ʪ��Ͼ5���i�E��0lļ�4��yi�B�Č3x)�ŝ�Ljx���և�Y2z��۟��$��67T�a-�����6����љ�;��;��C�����6yVJ����x-��B���@��jwi�z(ҡQƗ/��+���&n[A��Wщ��U\48�?=���:Wy��`8D�<�G�rL� ��mB֢.k6�Osx�W�����1�d��N���bK Ux�p߉��`d�Q#�&���͗�r����0a)��^R�Z,[s�R#Z̼��̜����s�L��E!��P��fH:�`�-��hF���:�q&��Qݧ�X^{���@!\HD-QN:Y�pË�=�>F�]�����'���z�o���yѷ(��0hy�#�2d��]�?K���}~n�S0>�^�&}�=��ͩ�¢]	[�9j�i�y������/G��̑�_�S�^_Q$J�b�?��J��D��`� ��VY9ї6x�ڙ��~w�2����%�f�EC*�)[֐�d�ғ�KSA��ssփ�*V��7c |�4Y���j��>�T�o�_CMv/���T3!���������d�����O"�/�|��z�H`��<�s�X������:�Y&�Q
��m%���%���j{.���)r�uW��W������b#W����Ҡ�9ݲW�䝌��#�Ƞ�^3g���>�!��$B���[.f�{NB['�$Q��&4����9�~�����Jf�B-����n��ި��z���LU^�(�0�3�MGM��|%�4��G*���[IK�%
���O'��5�����h�x}U�p�<Qsށ�i�=��~[������B��<-x�#N���2�	Tq�Ķw��Ti�_��z9�Y���U���ؽh�0��Q8i�j!�1�^��o��R �E��a�s��$iSm���g��oӺ������$'�o�o?�9��Id�Q�&���Z����i��*�zZm��f���U�O��H'�t}O�Z.'��5+*�jO��yE�A6�7^>�ʗ߰d\YM��zD��K�=:�K�����
�
�)8��dysAmP�����[nanA��ZJ	�����O�����F�ߺ��GB�XF�ͨja��@��+����Wg�B�ns����Z[��$+9{�d�G�d}�0�,2<�*�CE곐"4A��@�N����9���J�\w�����"�a���oi��L.�j�x �qI���̔i ������ھͮ���j��<��e���$9t&�����������?GD�6�D��0�2R]~�W ��.�ʺ�����������Yg�Et�el�r�$b��M��+ܡBS-�xmq���c��`��^Ԙ)ۯ���cH����̭�[?P\%x��i�=!���8m��Ė!PT���W�p���_/Z]����U���+8��m�<J}<؜�4<τ 5���Q�b�-��(�Z��R��H���\�Hf���d�V�T�����W�ca]J���;I�'Ӿ>���۷�v���ԕ�i��s��Bf�yƖ�<.�|��L8y[���\�M���pY��8�iL����~\_}T�p�%&Ap�Qs�K�2��/��ߔ�!�s�#n������w^&/:�hKO�6j�g؃͏����OhH����]��c�v��X�~{m�-$l�k[Jo�� ���8{� 䀵,c�E�p�M��˱r����5њ8A��0��>�tv�uԸ$��iDI�/���)�<oB����J��m�rj&�鎱�X�t���N���1,�4jpʋ@���(��/���V'��d����Tc	���-����ѧ8�/f�D/8�և��\r���A�{��I��1q#W���_�c�Ӽ�-'��ݚ����:L��}�0U��`���Ƕ���u���L
IYM���Q�8�/2�!�m���!Dr���v���kw�R��#Rtp�F̫˴"I���0�2��7�e�C{{k�!A��<��W�P7E�v����Y�u9Z��X���z5�ӬP�r�?α���,e�8��+���@z0����+�E��;f�B��NC����a��[�ϡ���O9�#i�v
��	,As�鞣��\N���2��q׬���!�a������30
=�/z\��$�Q��{��I����yt6�bk��1�����x�	�6��������<:r�P�uUS�$�=6"�9,��P����@�idOtY�bwt�aeB����]�l�����n�vj5,-�.�rV��|���I��a���C�j�R1�e����|:�~Gʬ]>�w �\���\��Mhb({|�����Ws[��l��9��WlI*��|8q���%�'�D�Ƭ}���]H(=���z#�yP�\ϛ�H�����WWH\�վ��1l���<e��l~2�N���|3��XI㽙�yFK��#��Q�Æ-����|�q��ȗ��j�Ș{HSki��]�Li$yt�#�V�+���=���t{_W�Ϲ<Q��Q��t}�8����xp���L[��Z1��#����b���IR�"�S���L�];��"�m�1�����ghӑC���S�1^�P�<R&T��dۇU�?];�3�/����e��e��X��bW����v�M��/c{Nm�C4��e���e��e�K��ɋ�3�����嫺�Fޔ`T�����Y���zZշ�.E��c\�W(�`f�7����;d`�ЕB�y��|k9	\	zEc��٥4X-�dbJ}��bJB�u|����_��]5�����4�\�[*�59�ª�	�O^��B}b~�4{�M�o�X7�g/�����/�Tt�=w�;���'���C	���K�1I	1/X)��d�
.��� ���,�ծ���>��d�/9N��
���ڼ�ԓ�(�,薰��7�V����.���x�
�}m)L��Zٺ�>:�w����ܳ�	G,W8��'�5�i�
���If�cd)`�P�iM���:9"��R~�	]��LL�*M���� 4-41��CIȕ�b����A=Hp�f�q 7Cy�B֙1æe�_\i�K������/�W�D�;�%ҰUS���H��˼(�������n��o��ڴJu>�01���V����N����D�h�$��Ln��l��~���V1��B��j�wܲm�f�WŶ��w~�g�S�|�Y���
��y��8{����RUt�@FD��Z?��N�e��������m<.c���g��ˤ��WS����*	cL�$��Θ���nyH�l��e���{|׶��<}��u@cZ�����(�54N�~Q��}H����N��ϛY�Í�h)B�*)�C�M��M����A��_M�V,={v�m*&6�=��35��D��B5*:�Y0�:�e�
��n-]����':����Ģ�~��'��T��e{YlY�*�������,��!��%�����߶��d���d�ΐ.��sYr1�j��w�^�=��Fҁ��8o6�&_�|��5���O��'������*����Y�3�W��Y�ػYw���E��N!Ȼ����CM{�ݚ3��M�uӘC|/f�_��T��x��/(�}�}b���EE���J �}���J���xܘǝ�v�"�����f�uw*vֿ��q�Q��'U�JW������x�"}[�Ց�ݙ�����
n�ܒۈ}t&��a��|���>N�n.���<��m�w��DE�9'<�ar�u�͛�4��VKn�ub�摉�%�.��`����g�I��v]�"�����ƞO�U�����~���Y�=}�&���gl��;��/�(.OPQb���"�'	ՠ�$�L�83X�n�� �}��1(/���Q�ū7ޛ�B��;�I�(�W�wt\���.|p�N0c.��o�3P��r�������NK������u����-�������Z�t�x����Sdt���]��@������X����%xYo����\%��Q�#�zY�+ �M	�0>�o��P6?��Ad�}ղ�P;/4=��`�e�#�¼<��,��ϖ>e~**a�$a�#�����@<\���.���-�&ijR�m��Q�`˦�j:+P&�����Q�\by���.�k����������;�,b�"1��ڸ@;�At�u���b'��|h�z�+n�]*%M����H���m���`�]y�����a���/��3�����s�_t!���
�:�3����1�� eOY�CK�3*@_��O�w����/Nz���"�j�+��y�؋�pk�����YtpcQu5���Y��5h��Ri�K�(��~F���q[E��J�Od*\9��B�����}���蓵<3{7e�Ϝ0?zT���L��{idg}un=S:
IOZ�G10h��b~���0x�;T�Y��6�e4a/�`����V��^����pu��h�wb��N!-�9tCj�
hYι�^��6�i���A�D��ѣFnRf��z�����
�<5�4kZc�wO-M�׉���w����"�eEN觨�m�	-�w�f����8� �i��h�y��vI9�.9���<T��t�QL'��E`�5���{��U��4�wc��6D�{m�b6۳�o�����2+����0����� A�hf�Z����
>�9"�]^m#����,��.PZ����o`�K05]�Elq.�+~����,�Ü����ߚ̀�W@)d�"(�[W���
����5_�'.��}8����
=�]!g��nk���H� l�-oB�Sht��I�*tL������j� ZEly��	���*Q�V�VM�Fڇ׮��\��R�t�'ezӢiy�Z�35 s�Ƀ���cD��:*�j��?V�g5L��9㶎�F��)���Pb)��t�Dw�H��@+�P� �O�3{#�)����X�����y�<W�l<�&���g'���h5m���d+�W�?���{-M�R|����/d�Oj�<#���
W��Lk����a�4�r��E=�y����3���r�hQ���LQ�絢bgRʠ6K'�GÒ����9��EA��������X��xS�U���"�9�E�QC���ُc%��7l,?#_:[}G�f�����}�Z<X�Y����/��点��?�s 6���FͶ��Z�2&Ku�������

-��W�C��E���ӟ���z2�UUp�݀@1����P������y����q��ʌŗ3�$����1���Q?
�{�mS�l����HȞ�5�|ŘN�'�p���[1����C;��c�;g�����k#�R�� ������q�Е�ǱS!ʉ���]H�M�P�۾�P����X'�ͪ��V=Q�W2Q���ͫ�����3&7��@	���Ԧ&a	���P�����,�LiuU�*����O@�v�c�&�Z��d�L��V�آr�$�:���j}��'Tc�洟���_��Z��]���j|t�l��.��M�?N����-S���MH�L��Y~��WWy����A ���7��b��VV�l#W�8�^�A0��Ј伀��N�?{F�k���
���^W������-N霑_14ވ���Ł�'�p���f�����W�i�q�f=VS��G���Û��Ltpw�w��&��=��TO�Ib�C�-��O��_�#N�A�/���`c�H����x��N���	���e0�����T˂�����<|W����2���g��Q��}��Δ0Uثi�4���L\�6tz��?k7l�����׳�JFt_�/{���Y��%t�} ^]�/&\vgj��?�����>3�`�dh�ΖF cǿ��rm�^��ɅE�va-*�7"J�E4�u;]%hs��>E�N��2:�eZ��rV@����$�fI�W|���������`���o�6�?Oσ4��K��+�H�u�+�~7�Un�F�_���G��g�w̬O}CK.��[d �����iG*��	�K��W~2 ���@�Y��I�=r!�� �c)��(d�Gx��d�]�K�щ��#����v�S�b�_�����=Ц&7��M�@��]-�E����Ȣ.�#�z~O���X�g}�s�S�w?/%�.�
Hۙ�i#rG���$/3��6S}��x��J�K���_�8�&�Z}�O�{��^O�/Oi$)�f6��jB��.;�^{E�w��7�x@*v���=�24h-Ɏ2[�q�=7-2L�Y�l
��tv5Q��?,��ff�J�ڠ+)��W� 4�d���2�������Ӝ�J8��u)��~mk,+��Y�����l�k[&�@�����E����g�Ph\M������8E�0��꫁F-��5�F�3�&"�_��G��q��f���<���H�/+�4u,=pu,<
�S�} .{BN������"I����;����M_����� #�#^�R���`ql�FP���m�E�x���irͳ�ʛ��y��UU�}9_�������:���6J���K�!Nm�=tN���Kf(������ī܂�;57����*~�s���sV�[�����2���Nk���&kZES��-��Z�E3+wԽ����Ee��%�o^�1��[�l�9Q�y���F,?�O濫*�y����Lɳ���I�|!jJ�w�o�I��4������~����3ۖ���Q�����QoYT􊩺�S{۵�nJfM�	���Lj��\Oˣc��մ�0�/��G�5�(�*�sїJ�ؽ_�ޣ��xMw���=�������DTJ��TP�����P�"�ѫO���6Y��Z|
�@��_����w��#�;k��u�	/��<QW�rI5��ʫ ����)�d:/����<X�qB��6{����9�K�����s_�Ӵ�7���Npww_��n�}qwKpw��,,p�������0S3�}IuUw�L��R�ၽi���g��h\}�v	��+B��9�˻F>�˟^�k���U�.��+?��nAގ�4O���uqY�д�)��OV<:�<]�9B`Fv[�Iʓa��&�X�-�x�� Ut"`W m#ë���q	w���W�"�h���K|X}M�hs�6�����^;�M�T<���̚ݯFo�V��GWU�������v2�r��"�<	:������a��Ҵ���R�~]7r+皰wE;���[Tl�U�vg����X�GO:))���c��L'��SS˂�u"BP��p^ڟk�9U_R�����s��;�s[t�;4��1��y���Yt7�C�ZJ\&(�J8Ӹ���\�	 ����1��k^1���Q-��%f]nkLJ��#����E� 8�e�S����.��w�A�\��2�PI��=�S�l�<�-+;{|@�j������#I�k�`�m��O�����4>��%M/o�f/%����x�/�3ַn�z�������4f�y�j
�&�>,�lo/����W�pb��q�]�
���PLM	�
6I�IIc��
 ����� #'2�����'�T_�����e�Q�ښ�p[�����V��9=�"���d�%;�M���/����V�K����\;*�Or�c
D��ڙ�)�`�ӵm��U+@Qիo�[��bA?tyQ���ԛ��ղ�{���o�9��eg�O��i/i,��j̡	諭Ɋ�[m��P_���"x��ef�jJT��Xģ��$Q4��t�ʭ�i��g���}z��y!�W/�3���K)�j�Udg�&z����g]���>��7n�J+	N�7
ҍ�2�_0ϐM�+�(U��U�<�$@+d)���\͟�3�ˈz
�-[pjg�L	��R^B�}+�������:���ii���U�5}P�1��JMأS��p��a3�x�����79�M9�=���Y����~ D�5��?�g�.�YScT�RV^2 ��Y�O��G�� 1�����Z����d�����q:Oe겦$���]zz�|t	"����9� ��u��O�١�����
n~�1��E��l�$S�Q5��Co|�b�\ј��Q�h�}�[�zve5��轕��P|�������)Ly??#Ёv孔��ϕ��%g��E�l};��-��?{�s<���F(Wg K��J��n`:�!sIdА�ֶV�N�ԣe�
������Go{��!�ϴ�$�[ \V��}_�pZ�211MW�?�Ay�M��X���:-��TX�7!�����LE��l!��F��(��R���t��>�d?�A�x�%-������#'Q�j�v��,9���Փו�Q6�d�a>�@l�LDڈT3dL{&�/�`����}�O%������ m��|g�7~|Ʉ�����ޣ���v��*��P��� ���s�B��q"�Y��S��	2����D��	m�޾��A�> �_�������s��������˩��6�<(����e\���,&C�_#�M�k�{��v'鿾x����l�)�tu��!����0���e����Pm�yez��Q�h�v�Ӝ��X=GP9-���V��`;�ȓqtI����:q��,��n�s��7N�k�s[1���V4���ӷS �����Ot)���˖�OuK��  Y@��[�6> nN����I���C��?�PG㪨�:���j�xJ��Su4��l[tJWՈٵu�x�Ȉ�$?�V�4"��q��z+���Tޣ�W�o�M �-����lL��W���S��D�$� ���n���ʆgo��ynC��krn�3�l!>>}%�h�QV]X�J���0���E��E�d� ��i�~��"ĦP������S�K�?��T��|'��v� �k�����&��L����~��^�+����Y�E�!`����ѿy�q��߇�채G�o&D��*N'�5��.&���'
o�a3��:���& �>W�-&�XH���UD�M#R d��.�4 �������r|Nh��=����9�C���� e��wZ�-�~�`ha����a�q)�� ��$�"�#?W���|�4�b�.�+.PPU�]D" 4��#���9~�1�9�͎.�ב�����P�gb詔1f�gr�H�@�S�� R�ܤ7�7"1��E�N�G'x�@�z���_�����M�Vn�o��)���U��T����2�A�u?!����9j1�()�߻Ϲ��Ѿ�"R�$$8�������|�����t�}�ti*f¼K���A\���,#:��\����'�B c�t^��~Yx8(8_�-��=4m��,�n�����?�8����.w�ߚ�����NB�^1R�ϛ�x��+V�����JD�������,k	I���������C���"/b�k�;����_�e/RG�ӎ 
(骑�~O�R��\Lm%ދ����UQ}�H�2wc�ȾLt�^�<l�}���z�n?�-W�[�?u)��2���%�/A��_i��f(!�֥%�K��ˍ�>]����^���n����A7�:���Rǚ��ߣ��o�H����k���XaÝ]��ݑ��/_�*�� ^���'B3$u1��(-".P���|o�� ���ljr���1��"�ׅb���q�Wt5V�2y�|*N������e%!���R�/��BV=�;�<ޮ3.�?^?P����O��ô�;v�D���ޓؠ���' �afj[�����')�6-�Ω��;�E����J�Vz(ت<e��P��Ÿ�b4t��$T+8fLQ.��l.#hftGO��r��<�M��ݜ�V���qF�Fɗ�0���ZU���|�R���3�44����'*�MG����Nq��'<f�@_��E䓕��0�<a@xk���gv��"A 20��㽘뽱%~K�O�h����zE`�{���;*X]M� Th��wF�3�WL�� �#��+t��;>��-�)yK���`���̱��
�����kmu�QJ�5����t�"�{�p��ʑ�& a�#%h��V�-J�K.睨K����B��ҩѯ��E|�l� e�&.ܭ�_�d�Έx],�xM�՝���{��.pUj�,vm3�e)Y<ޝ� IP��V�/�חq����_5�Bu���q�$BDP��^a!+��������AᥫJiJ]A2	��GC^��J^,���*AWz��6˨)��R��ٴ��i�_M3ҋ�)~�FS��Oʑ���J�������d��`��g�B��W7��n��[H^��Ӓ�j�'<���MV���@f&�H��z�h[8�s,���F��n�#&�1��u|��N�ɔ�9���k11�Rͽ��Y����խ>���v娇���g�yn1sX]!��
�����l�{{��D��3t/ߊ�&���y�y�D��#���v����20>Ҟ���$�����T��|k���,�%�*W6ȝ���*	�⾝��1���h�r��'YxJؕQ;�kR�P1�zV%D�|�L����	���a�J���<Ԛtx=�.�<:a4yQ�pt�D�&$ӛ&x�q��c���J̯"��.5�Le!��E�������3���cO.N���/�������G����tUzo�g��R�U�Q��y{	�����D�
a�{%-JT�ʴ7<�u���.��b�2��u��x}��"��nw��HPr�5^?Z�jlⱥy�0m�Ȃ���
�c�\��B9\'<�~Q��Q� �PR\Ă�׫s��G�b���\|��co��>����E�>u��Bc��� J�fs���7�2�ja� �K��R�Yr����������>6b���I�+,�+�]*��	�$�����9(*�JOP�vڱ#c���{�麯
�R�S+8^.�a=�����T*F"F��ه��4,�����	F��l}��g�V�_���&�+�7��0�ʱ���VV,�����4?�U$"�8A[�����y%C�6w�{6i��#������Z!��b{ߤ�Ҷ`���|%"w�? ��@����Lp�q�J;���_W�Z�3C%f-ijFf9�[�N��x��<��x�N��ФK~�hM��c5.z}h�{�q�����@�3؇UVb��њ�⒦��u9eq.�aٸ������򛻼�o�d��B	1Ã�S��~�'�k�K��Bck������13�S��Ǘ�;=�]ǰ!)�L=��%c˪"�5B��LJ��l�	���Ek��'m�Y��ĴrT1�2�w�#}١V���{a��'�:K�I~ׇ�f4��
�tF��!4B�`lM?��(,J�� ��爾*�~�t2� ���6_^Wp���!������3�7��ꛁ�͓�'�-��:�DC��t!nrPu��_�8el���A���V�DSL0�/�w�8��1��"�p��SOy��20�و�mHE2l��	_�,�V�`DM}v�����a!�'�t�B-��t)�mnr9�[#��v����H�Yp������>��^V��������7�j�3v�p�Cԙ��|9���X�W�`Z�� �(��p���"�J����q"W<r��z�X�N�L�S��UF�7��qC�#��ڎJ ��D(p-�/( ���q)P%��Q�)�Qzc�N\��a^�.�$Z��f��Nf�8��\[�F��h��,gB^��*˅���[��m��k�=�P.+�|��ڨS�@s8�S%��\V�En1������m� �K(�O�˿��? ��i�R������6L>V��(a�ƌ�ŭ���EG���G��;�JÀ�@b�K_�, ��򀰡�*�9#�;�Iҥ"eiy����zه��~ Ķ��N/�UV1h�i7	��5��������cEX�u$d"׵4���L����5�˨�����/ڌBm6�����*�-P���՘��~N�#"��j�u俕�?E#Iy��y��7^g[D|�2�*@T��~!X=��3=����n�#o_ml�؍2��yIT���yD���VNV�e9��Ǌ������ZM\��f���t�<5�%>��`�a��u�{�\��橩�������3�&p���L�^Ci�L����jvnZٻ2����6|�rz��dbˊ�V����#��G�o���ԛ(׽�9?�ſ� 9W'��a6��(Jb�vG*�߲7�V�����8'��~䣩�RhR��j���-E�������������IF���j�� �XτJN���=��O�5��$�(����쓧�"0+qI|u#�]�ٜ�"Zx�~���c�ǜ�j��� (��у��{㤧=�w��[!�b`�����t� ��.��.
�lW^��� ���c�=���`9�rIF�A�š�W���Sz[�Y��W˧'��(~�	Ɏ�n�rpw9lvP4�7�$��-B!%!T�1S���D��I���mͬ�=e��/7<�X?�g玘��ĵpR�RBz��E�H���o�샆SM�RL�~l-C|�zQ�B�ky�&� b���\tY\�Y��LA�ȷ@D%1!U���Kݝ����&̚���#Iɴ�h�xx�\�񩺼��nd�5-�Tg[�s�T��T�L�fy�3���G�b�1�^E��8��t�`!��ʫP����)5˂����AKti����3��imk�v|zkJ����x`�,G�n�x�'.|;8��$N��n��%�;�5��,9!��`�Ш!'�d\T5	���p[�N�C�EL�m��U@^��~Hy(9���0)���j�������P{������C��ذO�c�O��RZ拔H�%�܌n�}~��I����s���+涮^�`֙D߀I���ӷО����W����ūBf��h���h�Q֊�1��n�`����~���^^�	�3w��������> [_xCuI"�ܥ���Z�of�%����״�x�j�������ހ #|�#�MC���M��`��~e�M'{�V���%�kX�Ayn� ^�~��~
.��.�1$�fw��g֜n�V���'m
'O�i���ʌ7���{�H<��A+�̏�QYo�t0�s��&F:�6�5�9�	�s�G[J�WH��:`SU����m���dMT��[��nO[c!��c���h�8Io)삢|��3٥ �E����:�M�&���;n��U�O��C9�!3�V�� l�dť$)���`Eg��_'͒��m�L����@��bD7`����ŝ /����N?n���u �4�D���Tq�8�	�{2��H���Mt`q�>R�GT �-$u"�Ux��iM�6�_�=��F��*��vH 
�٘34W��c��fkT?�G.��>��m��Ҿ�C�<�$����aq���7Y�+gB�p&b�<p���Y�xj<H�gJ�o�:�eP����M��L&e ���%X�(f��j����C9j�Z�쐓�H&3��wTo�)�U:+��{���ԯ{��)� ܕ��n0�W� ��t�v���3]��@/����ʗრ�T�.�����lhaS�O�^?����&o5~T�a�&[&�'�˦�����!�,�| �����9��.~ �L -�o)��S�~M{����r�[Ѥq��*���eRqMr*D�U��I�$���a���F��=J��J�d�� ��� bZ��."�I?��qJ�[�%�q���m���;\U�e��m��n�S��\"�x{�ޖϷ���4?�xLb\� ����nC�a�֫��x6<6g����N[�U��ST��'ә]���;sD�0��P7-i����_���S�/�xWkg����]���N:�j�6��� uN��9*�l�W5�Q�l��9��n#��C���p)0����u�LΈ��bL�V �C`� ׻N ��U~�kDAp��������ㆰ���g���jܬ���$*FACg�8��ݙ�����VuݓFb�1�N=�ܿ����^�����Z��E���`�V�Ѡ��o�(����G:w�;����d�2��
lݭ�pF�V�g��c��B^�(�~��_�*+u�2AE�r�r���� E~Nl� 9`Q1]��z��ƍ�_z�{0�s�qY]N���,i��J'Y����o�3S8݊�֜^2zs�8�V������(ܮȋ�%�y�%���QZ\���&�w��#���;s0�r�9&T|i=V`Q���Fk��r����*��/x�0�Է��U�e�{�}M@�v�s���4�2�ۥ(/��uԶI곭|J|�-\B�d��C~�� �����{�,�{�چ��?���*ji��?;���m7�4{�@ʨ:�<n�@�!�� ��roͧW;Ijxs���'���kD}j�E��� tSOuCO��P��J��U�����Kʡ�ޗUn��u��!v��[�r��ֿ�3*�n^Y�����O�	#��٭`�ߠ��۹��[h��-���Ŵ��Y%�Fm�z.1�����*�9�TF2��x���1
�T��R��Dt��u��lzo�>>ܬ���K�WS\�����;�� ����y߽\�6EB�4����G_AqOG�7��w�]Z�5ZR�k��ॆ�B�u&o�7&�D<���̈Y��J���?�;��ka�(�^Q��dQxcĺ^ոº>��__�X���̕�����d5@I��h����&B�(P�w���� ��~�K���O��_t����3���ߔ:�7'q��1qI��.~;���J-[T�δ�X�aܫ�a�Ya����i�'OoN�ƿ݁l�-�VÐVǮ�WwG\J�4�f��'gʉ�V�z\�ܰuy˟;3[��U�6K���/GE#�r�-�R�زKH�z~J���8\i�x�!j'��Z�k�9\�tjM��_�kc$��D ��=����̏�SJKP�<����ȯ�Y�� $]�;U�I�߽�ڗ���j�a���	������	Eȏ*�I����m�g�0�$����覮�������Iz���_r�������p޾�/��� ~} �ޟS���_&V<[�.{�W��2\/�3��Ϧ������W��o����9:O,ʾ�0..*��`����q&b�u�<6����*��"Z.Z�"4�u��&�I�&�>���W�♧vn��h��Q鮽g u{c���m#�N�i5:�V����Mc��$nb����g� �"�]��XH4C�Hu��دʏ�C��甁sVn9��ˇ�ˎ�N���
��bX��&r͘�z\f������E���-�
���)_�ؽ�'���Q$ӯ[�?�dF)'��+TT�-(1} <�Z���ٝsR\���̶e��ڠ�²d�]룧;�����6*"���4��@�S�!��k5;��L���3�&��D���Bq�Onߌ�8���g�s��䃑���M�?��*0"�~r���{1F*�`diazѬʗ��%SC�o��#��Jj��U�{�IBb�-v�N�d�P��--_O��l�4ͯ�x��8��@*��"����p51�S\��gX����pQvg[�8�Nw����<��D����%����t�\"]���;�%��SΔJYOjr|w�b�skn��P���v��P����P��O;2������?�]j$f�6��0�%��6Usc׫H�P�/Z�s�诱ׯt���'iK'�������6bU>~ �<���M�"�=E ��0�Q
L�EZم����dR�^�k?H�.��p�#3�M ʦ4#��bc���˝íR���7c�*� 0���t�\N-��9LŴ����b3�����/XN,�KF�?�Ơ9*�i-%֗7�BE��E9_:�A�"X��ǋu�*�&��gخ N����'܍�K��u�`�K���ޮ�}z�����.�����ڭ;� ,:���D%�ے~����������o�g8B� ���>���k�˺��+�5��sI�((��l�2W$Tl8�/I1�{��N�ϔ7��o�xQNU�?�;�*v+��4@���~QX|��ch8�h��73��f��$,m�}�%�[�B0\{ʟ3O3�����ztn=��93�$h����/�Y#j�5Q��y�8x�(���h���a��u;I�䍥��.����>���$���w�� )w��p��c��%~�"�?�sd�
�U��uz*!��O!%�+K���">��+�g��f�C<�/�c�����"�ٷ�<���1n��XI�l��T�9,���F>#��i�A��Xtl�i��hAږ�����rwޗ�Sk�ۂ�hb�6D����M�~|��N���X������F%���I��z�G�Hɫ��h���� �p?���ϩK�R:���;��Pt/�n�c���u��=h
:S�tDwqv�˒cޱ�o_������yu�&����q'���)meuQ��{j�bi�z1Kyo~	��k�΢_�ؠ/����`�]�!�GFL2�C�5�cUH�2���3o�����删�׾+=��[
�����1��h���B�ġ��ٯw���=(N��Y�k	 ���0i�M��`
�^^DEEYJũ,g���]�9�O�> l=C�]����rB^'�E�6[ܵ�#�s�_�k3�גvp���s��G�~�(Fu�W/�{)�S�HHr����4��f8���	���`Z��A̖6Q�k��3��<���8߼�'������*j'�/&�j%,��R��:P�5������>�+����}�� y���ް��~�S�őK��&v���U~��EA������
^����HK;�d}�ļt�y[���n|��:���� �6h]��`�I͉��L������$+���~T2v�8%lj骚�2`ᯆp�؞;8ey^21O���')\��"4<�@q5V��ei�����)�824�O��o�ܮ�� h_��u�~"*ch�Ru8=co��P��W4��z�U4>��F���9����j.��C-��}D����L�3����u��ߗc��Պ����☟Ѕ`v�.�/?9&��4��xxM|�Y��sb�I@k,��ߝ&��t�lFb?=N\+��y�u�D�_ oM�t<n;/�<E���8��T���R�&΅��f�Y��vF�}�3�V�������31��H{���4�g3���hn�q&��
-@���}@BL�+���C����������F�|�$-�j� �G��}O8����	��Z���P��P?��N�Լ���S����g,��M�ˉ�IgDPݜH>9;��X/S&�sJ��R �Bz~^��J;��DB'��Eg�oY)�\%K����[���,ԋ�N=ҝ��!�e��4$���wc��rW��|�9g|�j���B�Ym'>�C��zD�K�S[�ЁW�TF�X�XO{WGv �C�>7o���`&�|�b
������I�qnx�����Y�n�}��pjÄы��z��c�!\j��=c�Lܗ�j�a���?�8饜���B���KvY\MX���L��O���6B�e>��/NҪ���Ʃ\ ��,0$�X�no��3��JW�!��%V��ެ��g�S�K� Z���	~h���s�n͓�N׷��1�׻�U�����}�@e�U+F{;[mv�ƥ�ߥC���z9�Z:���8�m���E��y���?��������s)�PmA��M��MFO���V�xb��N�@m֏�Ua���g�A���@�b��t�Cjc�TzM\ܧt��8�9�	�E�
<�ŵ0��L�ޛp������^X�/T1X%�dHʬN��p)`��đ�W�wR�/��	����Nj���[���	�ݓ�̪���O���,�\���;�u����Ѓ�%=��
M�G	���eZEӪf"�C�ÿj �MU��wU�S���ZVG�;�h���Y߿��C0D�ֺ������||���̆��{N������:�VJ ���.�M&�onM�Q}J Fh�x��ҏS�La��fy>��XCv/���CBa�Y�٤������PD��;�K�p$љ3�<=��=��9�d�����o8,ъK��E"�Egh#&t��YH8j�6Y8JE��1.����]�|���4/���w0T��fr�}i����R��t�I�#>^�v���_'`���t�/���,F׏3߸�B�.}ϼ9�}��|�7�M�kP�b�?z>�f�I��+6m�>O�����0����aa_����)�nJ�L�@�����2QX�/B!ח�2j���9�A�*+���s�@v�Jc��)o$�M{"l�P����|t��Y�hψ2��aL'mHG]���^�(�X��0��H��LM�L��Q����+Y Fk����kf\�4B�V�}�A��9��CMKK� �v�c��e�S���DR�^(��y��	�gMd��+y������D�/�N��S��'e�Ns�6-^^9�A�^#C���<y�[�3V��6t�Xs��^�*����{e}VI�u�E@41�p�F<�h+!��>c�}��.�`�~��z�9ӄ���nB˚��K���_�K^�&��O@޽!9~[(�&9\�����Y�ڳdg�y+4�P($�}D��_���p�/At��un�7k�!�1iQX\˄�������U�3�΀[K*&����@��5��KW��#8������y��Qs�&�)S*�� �e��I����	�W����+����M��L����M��_����:�%��!`+����Nk�����p��c�_$*�U]:��}x5�}@d�#�i�4N�* U�ͨ8V�=<\�AzS�V=����<�}ptE����R�e	�"Ðe|s�Ry�Nر+e`�������]ŕD��ό��AB����I�K~7
5�[Ц3�~���b2���z�N9¦!l�I��lyXZ��j<~�| R�1�u���t�ٽ����s�h��+��} p�sjm���֘��	�eggx줣��!��~��,r/s�E���fdY��׈��%�w�>5�?�d>��EI�$H��f��)�IF���ޑ�I�3�A�G����|�E�`�R�����UF����x.��v�t�':i�}u0u)Rz)���]�J?�Jx�4k�:�ZlЂ-�g|O�E��ŘN�C��a4m��z�0�+絼.��L"^~I�\��`���l�z<m��&w�B b����fG�"/�V~y`\�=k��Ju�b���� U�w��b�E^/�&��
�n��	E�#�w�+�v�6~VdX��C�۳H�E�p%��s&�p�b� W�)�>�"F�e�"�d�2m���X��V��aְj�g}{j��Vi�9{6�l��z���ZԪ�Z߸���B�;��oi���Z���3�F��i�/�&�ޛ�����>�#��V�M8��D�Y�����֤4�
�f<�R�_�~��xE�iw���2�a��s�A�-�m�������r���ܯތ��,���Źj��d�壪Ȯg�,����=GtgyԨ�ߑX�ck&���...��Ĵ��=%:�z�2��ucQ�jmt�����ls3��qd	�Vt
�Q�j�n{&c{���j�Q�׃��܍~%��1]Z��n3Ӕ.��1�����xz:q�l�r��U�����A��KE�z',�{*o瘃u�N *a���Ȏ�Y���V��ȕ	k]
�<�[���e%�����w��E�Z���{hT�G$dʽ3$΍�:<U͕Ȭ�x
DL����G��t�]7|��fP�+���GݕfWA�.X5�h��n7)5��ʤ��tm��˃g�Q"	N�n�zD�����T�?nG�dV��HNP�V�7*��}�鈥٪�؉3�:a�a������0�T�G���]ʖKm%���R]ޣ� �Pa�r	�(���M��B.:�`����$s�}G�e��1��d�+a����,�n�Հ��m)�qD<�>rS-����f����е6�9X�p_���z��1hMy��n��_��%r�Źg׊���U�f/ur��ß�<0Y:�JgtJD�vT�5��%�P-rY��K#t�I]���/w`a��_��>����}˕� h.Qm�$tj�K���Y���w�Y�ja��/H��bϮ�wz���z�A	/�Sn�]�,F� h��3Řr�����~ ���/|)��r�K2�CU�? �U*������|'/\�u7:��f���Z`���㓲�I�r~)Iy��.��Ɇx��x��j�
c_����0���?D|��LG�Xo:�ް��F��#x���Ѯ���q���T	���jcE�5�_�{VMc������-��vgƌ:g�&W0��0a�R��F]�4����Οg����h���K��n�>��ϖC��z��5�!���K%�8�@@���t�V �sG��|�
-� kn�5>>N��x���]ol�;/�/�1�!�z����K��1|�z��;t�Hs����a�«$K����0Q���e�x"��#ͫ�(kRBV~3��!��'C'`zXI..l<r<�y���"�{SX�[�#~ZX4A�d$`��t�J�Aw�
oWy��/E�+��Q8���:��=E���W�&�o�ۀg8��>���66��`�W�y'C5�]��$���w���!�^懖��ɲ��U��O�����p`@�yp0�΁�*+L:ddx fʟ����R�<
 ˴R��}�8�%�Vtd���Q7y\Ċ4@E{��|�t+m��³�#54�lr)m�L���	WY˷�vY�f��b1&�θ� �iN���`��}�y����I>�:���g�*����� ��b�[
_:+(�(U�$5�d]�5��Jq�Ty
�T�)9qRQ��#����J�
 EK�]1Ʊ���owR�<�)	>d9�HK��;���վQ��(z�U�ڼ+"��pC���Q�]2��Ɛ��b*���f�a&K��&�e�\���tS�����d��w���'\��v6q�FE=<��(]v�%�h���|㪑�{���Ѓ7o���ԛi�6�᭖UP��M��	=z���F����*!\,�9�L��--�i.M�1�j���O�E��G�������T1~�*9�����خ I�p��W��[���D��"6���e��^M����n ��o��.!�&�"�HZ�凑GA'���.��w�����6M�����s���@(@���t8`���G����|��4���fk痁�9}��ڂ��N����M��k����!�K�X���rgY��X.����)��io�A��`5&`_U��~MP�!�m���l���Q�l��Z(*ƎҲ�����vc����a�E�=>�M�t�4�s�
yd߂�r1�~M�,ΡT��h�5$�#���Ȍ�� my�]���2��I���TJ�Jˇ�)�ٝ�~{Ĵ�q�$;�x�s�aӊ�R�Ec$�:�q��~�s�K�'zW��}|��ڢ^#�h&?g����4L�G����T��,���hE�.�u(�a�=����07gź�����1��8�|�Qg-�o��̠�؏� ������C{{x�C����sCcO%�����6c���\mj��&���ٙ��L�9(���o�:d�=�#�Bsϖ���~�MNj�i͙+��6_�'(]qU�F�'��H�Y�s���E�a�p�� �֌B�ڂ�e�_L�\�ft
����f܆3E�/����s�$F�;�ݟ��8$�N�@��T�<=�Ol����$A�w ~5����O ����������Q������NFQ.��� ���������Urш&�r��^����q�[�:��Wn�m�� ��T�no#�޳� �:���f��71k0!��.�TRQ�[r�1/=���/�wP.�l8��jv�}՝>Ϝ�TH��, 1TQ�eQ(=M���)����U!v�(�H�nD�:���@_ �h;i0xɠ�xu-TT�ǣOT��#U�ڲ'���2��i,.��`�r�v��"]28T]2WZ!ڋ	
`N�eˏO�.��7�}���*K�@�S���<�(�k�+�^�}ճ��Nܰ�S������5�#��#�#��h}�V��~-%���z��m]��c�-F�n��E�$2� דڳ���^�D9�?�A�j����l���3Q�����+!��3��S����/}�T�6���Y�Q��"2^�O�G�i�I8��_�i"=�ް�tG`�ފ��3����XY�@��̠"�r԰��R��)��V���W��G�_��h����Un��I��h��Q�ڪ���m+������S5�Tͣs�t-����~u)�������W�.5�(��/S��&^w�J��6�i�/WpE���ª�Y,��}�ְ[c� ],E0S�}	6��,�&���S3���i�©:|��=����)���h���k�܋F�d@������E���i���l�|և�Qyȿ[z֙'�����#�h�7���q���xSa�\[�r�U=ꄾ�i�3���#�<9:;\n�R���#\�#����$���e�,����@$���i
�ݱU�Ћ7Z�1�����'��оMX�+���5�?�u��ߋ9�)�0��"�!��r-������o[�q�R�,ZD.[D���"�O&M@��h�	�q���P��9�sYJT����+���!WRGf���e&�i�$Lpn�d;e�v�h�d��K`)^</O��*eBb��0��$��6��Bύ3!�&@��>�2w'��N(mR�S��|Zx�=��\`�����������3E���B1��U�V�%!&w��Ύ<�"�N�TMu]R��	�L�m4�-�@5S��N��k�#-��`��F�x4I"'*���y��ʖ�$m�Rg,�1�����^�G�؂=U��yx�1m_��|��R����ڲw�ٔ�h���K����(}�Wm��[2������n��HI�J)9�p�����BE��B����oY\�Z}<=b|2�4m�-q���*�xh0�$�mr֧�|=0D��#iA�b�
���,n7��YCmnaQ=g�-�
1��#U��޿-|]��t_B+��;\��Yh�bZ[�ly�
d�c��K� �>����M���iR��c���7����� \�����93Q���>X:]x��|��K��f�_wa��l������A�FP3c��b�㻽S�CV���>�NZ��1�Y��XaQͩ{xq��0R5�O��R��ڴ�y��<[ܗ��'�ة��F@�k�)41�:�V�O��w��34DѬ�����|�	�?�N8'݁��&t���93�?���-
7X�+()%�H����Kww�4��tw(��t7Hw7KHK7������}����3s�}_3�Lv{WG�����Pʄ3����.zw�Z�^M-Շ7�}��f��s�ƶY.��͙����}v��w�hˇ���jנS�5�����������Kn*�?�-��լ��� ��I�c�l����Xf2 �J�|<ܴ�9�gB�ùy���P���[�S{�T����R6���(E����f��b|��_�c�cϞTT�w�t��n��ȦD� �%��#ܧ(��0�N�/�)�X��'B�������*��� s�"�t��X\%a��}q���/T�j�P�p�h5za�l�x��N<��j4~��u���V/J��*��4����ur�vo:<ȸ����kӽV�k�-e�:-�{�PuZ�_�Wo$��k� "<x�S_��U�l&�0ut>�Vs{�K+�EP���> -��,����.	��������ӭ9GY�)x���kb�J��i�*�����^K�}��( �G��ߡ�kO��|[7o��?�A���S���6���u��q��bC�@l	��5dlFS�k�J�GO�-���!�5��D�ڌg�=�f?S�]�On������r�*��w�K���٭���J�MK�����_'��aNݾ8�e�U�����Я/����Y�d����ۍv-���lr�̐$r��<�*�'+����}����%��E�x�p��aS�Q__\A��з�g�V�8��[�*�Z�+��*�֏bؾex��8;�`�
���^[	P�Hl�ߤj���o�'�6>��#�?��E?��� TW0�>�F*�J6���!;Ql���o~q��߫�=����4�����SQ����.��Ntͭ�P�h&~��;dE���x��w*v��[�OG(��B�v���dP`���?��yNO+�%< �91+%���a+�k"�X�QmbS_�߮u�j�"
��i�\Rw���A��d��̭m�JGT�����k}6�?Xc�xKX�0?}�`���=�W�@v"گ�M-�Z��T�c,�����Sza��a�{.gպ4�K	5A�/<'jqb�����!JŲk&�4���q�@�����ڧ"�!U[���M���q]��|㴟(�A����;�"��I�9�f��o١PN$`��=�o2o@c>u��ږ��XC��:��:q��O/Rއ�t��4H�݆�+��|����倩�Ա	U�����{�X��ddԚ�zvO��c�ė|+S���6��}e��)�����i���Ob�! ,�����m�����ʬ0Of�\�����$�k��BL4���I�E$&�_(e�Q3pQq3
K��Z�}I�<��x��0�_<��a�ę;�-���ͫd��ʝ���|��/��I�����/ʚ�6:R�Z�n�����`�Z˞��0����0
�x��UsF�
��d~;I�j/�'\��֥_MN��B��W��0�;ȋ�F�QĂ���!+��I����_�S�e�gD38�o�'�(m5s�o�O;�~����p����'�
!��kTfVi��i��if�L޼��������M��X_h#dIB&TW���MIkp�ǅ�w���Hir@�#���r�X���r��g�&D�u_��QYr�uW�""kvw.`g�jcu����f��ͳ��Yɫ�81{�5y�~��nz����,|J#�E�`'��"==v�o7:���&�%P@�g�d1W�M67^�s	Q�O�z�N �ws���d�|b`�H�8s��O̀�2�0�<��W
�1N�'�ӯ�.�v4Yv�����^��GE��{~i�Ψ3���<�1p(XG�(y_#�����Hc�DSZ�%��nγw���Zhsj��j�;3��h*)rR}���Y&�s��������}��1�w���b�� n2㨈�@��'� Q�J�-�6�</�kjkJ3*Qx�I�Eb�m	�Y�uՅi�2f6�CM+MF�G؉HK-j+s��6�*vY���%�&�ԉ>a�m
adF��r��_��Uu�Z�9�u�aa��6���� B5��k5�:�X��Î� x荦�=*줻�_O��m���k��{�nw�8����N��$m���3�N���N��ZC�B�8�<=���#p�����DHh1��Fă9��ݽ���c�,��MԻ[��J��c�_����s��ӑ�&P�ԸZ��D<�$��=��%6~z�_a�r�K��u!+*K���jC�� �d�MY���������֥1��'���q��@%�U'�SX���{k�L��F�����҆A��7�@�ñR�`�E6z��	�v֒��~�_M�s�J��Dc�1I����Aw�L�d� A�R͓���+�~��H�Y�^b���	6F��K���3�M2`������������׬���&7�ʳ��w'�]�Kx�f4���4��?�vf����0]Q�v-nqֳ��Z�᥵�JnI�
	X��x��y���b)^��5p�W ?��~It2���������;O!.�b�\tuU�N'�����ʅ�Ae
�gh��=]66&T�����87�㛤g��$寀���^C)��p�����p�Qn�*?�t9�V���^���(F?�;�V�°^�ff���lYقLeΡ�r88�H����$�3b�JX�ӥ��}~ �7�z�J���ע�a�Ȋ2�O�Xf��m��G[lvK��
�֝��z~��,�m�j-RhY�W�m6�Cqi�8�ԋ	k?ޯ�Ο#g'{�zw/�>i	�b"��u�d��hkU))�qS�3_�;m����#s��`�Ũ�����4觢�H�.;�)+haz��.��'�|�����f���8E�����$u`�������h�Aӫ�;=,�J5$j�ޭ,��y@S�!����rO<Qd���� ��?�ϔ���@�'���)�`�a:�sX�	ix���-s�#K���`�,E��l��g�!n�fafIͨ#�^�fGCc]WL3������~�O�&�tq��{����)�<����ƒW�ѬE�tm��.��%��+�ȵ��ܓϙ��mlp�@mY�-�2�y��}6��L�?62^�K]��פͫ����2�O�J���S���/曶��_4�\BE�1C��%G^�+P���Z��t;��#���I_hi��D}h����fI���H��_.��&��8��_$z�nzo�	ܹ UoU��7���E�������U;�l���%��S��Z&��	�v���Aa�m�ݖ2���4��Kjq\���U���@e3ӊg��a6��?jߩ�����o�OЖ6hD¬L��g���Y��rTkL�[1�I�uP�NR�M`�a�ܪv����2ukp0��'��N_��*Zl�8N7oc����-��r1��u��_��`|������:���:���.TVn��������ۅ+���U��"9r@E�R�N�ҽ���<�zĶ��9�v���W�Y��vW.�f.�𳗑���W��s�I�u��hf_�+������5�p�E؛�����Y�|�V-���~pz}�n�3�|�M���]�D����N��bI�h(�݌���RyrXtz����hʙ
3A3�J���J(�.��=XRd^ G)��1$}������J��;�3�
��\�&���Ə{s<�
H�qzpl�^�l���ؓ`9�A#k���3���NN��BG�賍�Qs7�s���vf#���ot���V�,
�i�ѳY�FѸ���Ҙ�����33�I��b�����,)N�Ӵ,��������c����r�Rv+��u�}Y�����a�ۈq��:�8e]N�Y��oI�aW����y*����ay�I���.�j�W�˖z�z\~} oa$�4Ӕg��]�A��	p?�[u�4!h�EH�Py�˭��@PF�����fK����]�����_�(b��&���c{$։L�����5��&���҈b$n� es)"l5j��'5�Dd�Iߝӯ��3�i��X����л���\�_���sR3��������0HN�Г�u	�\��G����"��\.hlad1��3���}�=J�Y�6. �?Ͼ$4m3O�9mH����X�r��;]�v�;��'����*UQ-��{����M��p)sD�:��_����s�|��MbV60�}���A"�P_cQ��B�76�D=���Zً�T�)������]ZZ<�=^�n���ݴ�@������$L�:IB�7�2��N����?YT�WȥH��G�(J��n�J?#��0��uJC�w�&OS~��$�K<|�M)���bg�MʩtJ,w�QU�'N�0 �W-?V#����"6��l.�nt"�+�.h�w�AyX1��&:x�ϓW��r���&�)å\>�u��>`Ǘ#g�,h�tU��$Z#�3�~Uu"����6�۽E1�0GO�TӉ���u�p����Me]�ګ�{z���G������Ģ�sNVĲ�T�$���L
2��2Wc����o�S��6��w��Y]��|m�7���+{��"��+Q<�;voc��(�x��554���)$�Y�]6=v҆2�?�������̗�P���m�IXl|�/_L�yr���,��d5�A�MX���9�4�|J��y5�*�0r�&j�1Y�X2�.vN�c�vY��t�"j<Xh;��z'8{����ه�M3e�'�v_-b��36Ռ��p����rט�Xhk[�f{Xҹ�!f�"�(yݓ<)a˿��
µ��pҐ���[ˡa��9��Y�1[���nl2�CZ�d}��~�I=H�P]�T%���|���w�#p=5I�p�\C(�K&o�ZF�z�Y���ܤ���B�7�͎냢_�/vJ�F�+ >)\R-��/}¼�p�0v��#ڀ剱����G���\�0M|��?F�``�z��Q��e�w� 䇹3����RQ�S6<JR�&B;)�$���U�%�b>�p��\jҡ���96�џ@YI�7G��p/Nv�9y:1�`�T��(*�tZ���.��G�眩t����/$��U��J�4����wFБ�'�e�<�k�9V�;���9�4t"F�t���: !�'/,h],ߎ�5!}����@|�@��' f���:���+��7z�y���>(n{wrh��w��|�^l䘙]$ʲRf|�� }���m�����.�.�.��<�?p��'o9�q1��L*��5>|[�{}�ޖ�MO���6,�6I!S[��p_M��J&XLK�*f��"��KQw�x�t����r�l����nR�H ��6��O ��H��ӂ�@�Q�W �ŋ�b�`�s��bb�`?�W5^H��i�MK*��G�65h{�����Ǌ����fl7�.w�s���o�W�3	�J�f�\��p��]���%C�?��;.�0�����ۨc,�NDjߧ)Ѿ��Tߡ>�i�p4hEe�@��-CD�?�.$����/x�����F�#T�r#�Ft�h{�Rb1-z�ߝ�Uv��w�pH7�z����	ş�6�/'QO��[�^���d{������
?w�Jk᯦!�E�Ӊ�}:h��^*˷���6X���-R�]����a�j��#;��ٕ/tX<���'=_*�*���&��Pw�8��m{��_���zS��z2t�5AV� F����Ì!�'՞��a>{K/޵3?�ҡ��Ɉ�߇6?�>1�XTU�8?�T��*�H�k��<$�?��[@��&a�W'���(u��ul��R,�^J� �ة ��@Bbn�e�X�ʎ	�W@��7�GkKD/c�D����ÈOH@�@�����j.=�'�;��w��T�����i��-�57��]1v�k�1�vKp԰�g�S���>�8���&X��g]Z5�rALN.�Ho�-�����X袀���P���e���Rׅ�'I�E��վboR�V:H�E�-�+��O���sfz�N���u������!�uwU��$9�=����.}����=M	��CE�j�;��d)�G�`����x}J��PC_Jvb�6��+ �0�Ҿ)�x-߬��	k:����Pq�칣�O�x���0aR��S����At���cv��k�kJ�F����j�(Âd�۰�F2r7�^5F黲�}E�'��O�N����H��:U_��;�OzvVq\,��CVԁ�K�ʉ�Kڠ<��4�-��P�A��c[�y-�]�9y�X����몴)O'�3k��b�F�6!+�\q60,_�B������u'��QR�� q]yƷxm"�Y�z�c����� Ŀ�Nf!�]o7���M8f�nl���4�A�m��s�H��y�O�zl�;�B�NB���/�������{>W;�o���`�3�ԙ�8��c�м��d�g�}ŉ�3QDc���g#����9��u��yǮ�UbH����{�jJ��[f�NՑ�pt�o"Z�u�t���O˺x�O�#��88���*�I�	�/.�='���iE�ʓF�tڛ����c���P(zm�����u��@R�N���&-�����q����>�:�{&6�㮳�����-��,[�­	�,�-� ��W���䛤��A�4^S�Ky��.��%�+���A���aH�N	$4�r��1&��g;�.ð.����V��b�s������t��� ��fn,�P���D�=��R�K��Ч��W ��	�K|"�}n@�N���P��/�*8N��7�F8~�~�����{v������-U�5��,+�$�e��/�{�u�n��g�2��f���<O���Ӓ��D<}��F���pF��zVM� �۫��Y06\�򔞶�wJ�"�V2����(�$�I�T�7��b!��S�Nc����_�=���aI�j&UTe7�q�ki��6zZ��n�T�Y���s�����,�"�� ���HF�5�����&Ҭ�
��e�1��*��
�JK т�Ã�%�fo�k��2��
�F�4T[J��P[v�A�����L��z�=K��7��iE)wT��y�j�߳�I����u3�l+�^j�E@2�i_-O�{��Vv,ߒ��9Hv��b�x''�1���K�=t4በ'�OC��	uh���+��0��g1١*�)��4f��y��i�k����C~��Y�D�S��G�Wz�đG��j���<��%EeeOmc>;���h����J3ۿP��������[ӷ�����q�Xi]�ò�X9�v�ui!$YZ�\��)B��a���g,,���-�e{i.1�`^A>=�KJ��]�/�߹RӰ��	)��g֝�V�D'҇��q���h��P%a�������� ���5)����JPHBr��S�.��4��ґ%���I���|x���y�ke�����(�ʋ�xl�rl�Bd5�\�fJ�|���������~��D��ݘ*J
-�$M*��=T��-N�پ�#�=�/�r�`���O�2�{�9Z��מ,wݢpl/�@(��b���hL����j�l�f�v���t�.R��I/Es+�>���/EϺ�](y�y�b}��K� �5�X��3����N��ˢ�,�����0,��u=8�kda�0*4���LF�VO_��)C$G�4�=̒�}�T��E����|��v���_YZK�mS���3���g�)G��8� >G��(��R'�쟗�e7���zf/K�xl�O�]=;�P��3P��㉯,�$�XA?��2�0]
E���ᬵ9�� ��m�+����uw��|eD͇!�.��Y��T^*�9dDT���K���ɛ�L���\؝��a\r{��+L�H�3ͽ�����Kym���ߛu�[?J�� 8CwZ������������5o�
.��N�*Np�һr����n����	�/���䐙�evm�*U����M՚f��ph���:(��]Ͳ���JX$��o�4���$	u��s�i3;@�r�D�.�]�K֕�=��:�K�O~�U�%�J��`�U�4}��1kE��`�[�at��\�Q�rFv��<k�J�i�bL�N5Ap��{��q��.�M��ڊB�+���/�9�imdFḣ�f��E+�*D��@�w2�{˦�kk�Y������*872��Fi+¦���ℤ3s�)����Ȱv�sjq�rTX�+f���Ys�<�|��v�_��-���E_�A���mF���c�Cd���]�����y⧎';z��l��oB'���'\1��i�M����#���#�t��.*<��3��ǎϣ��#�r~g�,�̺흻�[�fY|����"`�.�&!��Q��F!�z��OzM!^�����1�l�o����:<	����t)�-��#]�
-bb�~H�I�s/�=e`����=�Y�㽘�<���Y�處�f�S����)r����cn���+`����a3�޾jB-��=�� ֳ�©�����";�����mz����D���� :@q9����Zm[�s�+���F��չ��t�]*u�����?���-m^ș/�q0X|őQ���n;JC��2�P��Q��<7��/as<D������~�������8�pó�G�j����7ǽ�G���|�A�^�o�#l��%縊y� ��n�5E�:��4����H߭d���g���A��ѽ8��춟��7`������pV�~3�Ǩ�$w����5��b8XIdҁ�#k����U}�N<e�5R��W��Ŋ��^�M%�}�ؖs�;�V]��KTb:�������%,03���<^1�OH�� �zm�V��vY�T�Y�yD&:q�|0޾u.��v�����N�n�V5$^s8��#��|�a�%�o�,*�y��&K���r�)R�
ca�LW����B���
)�M�9�]�,Ԗ�#}itlX\��eq���*(C�}D���:tJ��o;���-����P�������_�+',&�D��܋�dmN���~y-�@hqH���|X���΀q�d}�\��P�e��}�rQF��bwdќlj����"��
�������]D��^[7Z���+4�.�sG����T�W@�� �9L"y\%$�K��SME}'�=U�[�����W@W�O7�u~�����
���'���C}��-�P�|�%}NlZ�U-CH���s�|Pe3Q�S���_S�Y���O�-KB,:�����6�[��}�f3"+��Lf��(K�4*{�\��'44Q��9߸�o�]G�X�匿>��<�R1��!y����q,j_��_�ܑ�t0�N�����mu�3R��t��v�r�?fzM-�C����yS��|O1�
���H�mu�ZަM�Ws��[�
��n�l|�+~ͥ[��� ��;n��Z8_#�%�o�vay��8�~6�o�����~U�L��(B���M�j���m����oV�U��KuM�M��$�8�}��y���k^IDoR����ܔ�7�S�R#=����ۈ�;�G4}]�sO�󈸭G��qd/H�����LI"��X��(�M�Z ����B4�>��f��3׵/��{)���M�9�8���Yn�<v����nb`�����z���2�3�g;����������H��V�X_U�
�{�+]ˤ&�B��C� ��];//R�]��ݥ)�O������{���p��cG��_ڃ	���х`��D]�)�	���wW��ss�0���#P�nD���<Dԇ��x=�h���c��8�����=��2ɾ��A�?���K_�>c�9^b�v�U���.���K�eQ���02ȮUW�8�@��F�t*%_;�Hu�HM���6��&n{�u�	���zb�-�ͳ(�I"(z���y�n.���"�6q�_�#�����W U�Q@ԆޯE����	a�Zjk�[�\�L���}�UT�%�����X�,�I��u���U�ʫ&�"ħ�6�;T��\���E��>�֜��D\��E����	_�Ϛ�ڷ�U՝�R2��w��]�w������ɠ���dZ�Q��#)�M1ã�n_o�`W�ȍ�T�eE���`X���Ԣ}5j"̶���������bvc��T����\���*&���n�nKd���ۏJ`�����q�uZ$qi��� i���h.R���1L$��h��쥛�S���U)5��w��W�q��?'�(�4>gY̘�X"їt_�E�L���1�pn�	�$��?����:�!j��yDb7~jH���A�DW��4���iX�sނn�*��	��?��cH��R�:J�T�C΅��}�P��k�cz�˲���1��%�m[M�~O�OG���=�.9:�aA��J]����Jʛ}��w�!����E�jQQ2au�X� ���c�Y��1�X��:���WTMG�#�)7�,zw�&1_�����'�0=��
h0�Z�WI�?F�����3��>o�f#���Y+{�g�Gw���{.!C�E��96V���Q؊�a\?�[{�i���ɻ��9�7�fD{��ZR<4#-M/�`�},�����%��UQ�8�k1�.P���|F����F�yT;��M�m�ػ����
c8��D���=���
7=%���\�Ag�]{Zy�ӎ~Lږ>P�G�L�:s�㥠�N�Jhhh�g*����i�`f^�-�2&�8�/wH3c^�9��IVvM��t�����P�&ɚӉ��-OE�{��p��|��m_�
�L�,�X�ȵ����,��r��D����. �F�z��r��h��7RWV*
D�}���=�t���^��49ʽ>�QD�L?mP�Fщ8�s���B��%K?b�dݜ��Y�΃��t7���Ʋ����^�L�?�8��r�2�r���+CM��@� ��x���&��������޽�r%Y��N��vC�mmO'�L�y*��I���um��>>��<r���f�����s�'��/jsʚ�_��'��.����#_��T�bꇤ��aʑ%�qz�L%��9�B׬PT�	����d�:������_�����l@�;+��������"�iY�HI�kGP�1�5�כc���m}O)H�K�w+�����AX�b(9�My}<jv*�0們?)vѐ���{�6Է_�N�������&�]��RK*UVb�o]|��whQ�����w�i�빒�q(�|�NC�坺�y�b��i���5׍�}�\�����wh��V0���ޕH���<&|3g��O)a���L�qbһ��?/mE�D-wB[R$w��5����(#hZ�#�(oF��&����ҕ����aC�H+:�y��Yྀn�����;J�1G˟'6y1MM��^yV��m��?���s��
����<��+Ih/��^�����^qG�rIdB�BhRi�
0|t���o5N��y�<��ɳ��jx=����R��V��-��7�<�!<�,���,��� VV�SG�=�J�z��g�<~��NN]f�k��g�`�vlE���r�@����}h��V!�����?p�'�fd�D�3�֍{�d\��"��Fo��,����7��3�=Y���3��hI�Y�\܇�1��\���0c�y�?���:�{s���F+����A�M ��h�6��I����Z��/���,AteOD�B�� O�#�\6b��'A���mk���r+?mK����^Pc�����щ�RMOO�b& �����<�+��e�>�U�5�«7�5x���~(H٦#�1�a��|�g���6$������ZjBl�E��|Y��_|yM�Y��t�?N��p Ћ��~R�!���D���-gVP �):�=�9;�jqs붿#\B�I����l5�x�M@> �M��ɶb���)�����ˁw�O!���<�(?�}�����[�#A���$�����x�ՔL	�jVu5�Қ	��+Ja��D��	��j��$�i2Wօ-�'�o�8sp���Q�s����Q=N���s�I[ٓ�T��ۗkhC�Y�EL������`CTJ��1�a�m�����z����:��z��Nو�/S��t��?(����4�	[0c�D-�atZS��F�{�<�sy�<:��MBR��������H� !�
��P�˱'�s,���rM�U�.��
�.k��QX����f�}�-� ��$i�%�� Hww.�k�En��vY�%��&x�K��a.�(xF9o��<"�:���U{0=�}���l��[̦��,��D��k�xm'�*�˫�������p�s��!�E�l
�b����Fv%v���z.�b<?`�PD�<�d�Y9���V�n{�hK_a�ʘ.o��eiA =�eʃS��.RP_��HW ��6�W��>�x\}�����+@�ёJ
+{%��UX��|��j�n�7�7_d��I�V��aMݔ�*
"]$���g�i�O��c�
������q{ҌyOHO����xzj6��Oʨ��"���v���d0TU�!�o��I�(ph��?��
�~�#d�K��cX&�[݄X�-~hC:uvt�m����1���s�dN
ذ�,ָZ��9i�O�ۃ�x���C�,\�RI?�S��sp]:J2���HF1�Q��C�c������M������e������C{�V_~���F��sﴛi���|8s�s |��s�����(]yc)m��������E|n����kb���KN��|�jʹ�Q�DM�d�ֻ�j4Ꝉ��{�D��!�bBC�x>���I���.XN�f�c��8�O�����8�C�����9(s&<(6�cX��;w���t�fBjE��(��$�U>�
k��S�a�Sʹf�d����67rPs����غ�_�Zʙ�e3��Ϡ�m>��,���)�D����H��y_W)z������ȄW��n�_���'k(~��R�u�h|�g��j'�^I|S�SVȆPX���i��\��s��E�l��\F0����eH��fq�[�9�k.AR�av���Lv��~�>?4|�W�R�]��$-�Ab�%����;�/��QX9; t�NBUm�?��uU'O�.IyN}���<�`�����ٝ<n�p�yݝ���щ�y���pϼ�Ԫ/��z�F{3��D��"n�Se$��*6΃~]�w���V�2��CF���3Z��ɪq�Kӵ��7�*P���G�8�A���5!�}1U��cM�+ o���Jæ^��J`����e����S[��hW/�r�R�Ի��d���]��ԮA�R��+��{�m<���� ��T�^���
@`�L� �_�j�W��rv��lQ���';�WD�"��^��f~�@����=�$s{I��f,7j�C��'9Q��|��.��)ͅm�:j�pd�%C-��{c=m�& �7�'K�w{���>PD4���n��\���<4���vr���=�z�V�歯�o��uvH�Պf%�#٘#;�+����_~z���(jcz�ॱ�9�/���itYR2���$�x�����D�
�{i�)�������_�����5Ҟ�f�;�¬�r����M��,VW�Wi|����zr���z3���X[�)�'����.�����-��3n��pD���+ �݋�m2x�����Qa�{����iu��Lvn���$}����"�`g����[b��\���i��#�U��Q����4 �(׏xx$iѫdۋ�/�N&O,t�w�D�HHbA|ku�w@4"֔����wQV&��=Mb�>�Z-��dbj�̗@Z�CF4NY\�^ܚ��n���+�:�t�����V�>���?�\��^�d4���؏����#��Y��ׇ��*,YR�Cy1!�1�SL���7��	��4���h'�+=z�:Q�_�z�85�2��F��S�����Y�{# pbĠ��|�{��5�we�h��y��k#�~>��P�?[gt
�>��1Ĳ*�F���:@��k�쭴������|2�&A��oU�rZ�)o���[32�B][�b��{�l1�����ӧ_Z\�B��-��G���;�e��8�tX����>;�+ "%�QFxᄂ&2�i̞$Q|�`dp�2(b�9�f|j��md0a?!C*���Z.��Q�h�h��y�c�1[ٺL	z�:�RV�D�UN�S='u�aBE�_�M4~�]����
?��,u��,v�ѩ{��oz(<��	���dQV�qe�;s�~�s;��"p<i�}Djw�,.'�*�,	�/�a��	��Y1b�y`�@�§ڶ:�����G2�ҭ�C�L��m��z��A���@�ѽ$��<m׊�m�ls}��U�ۑ5�,�Ě��h��D��K�N�O�<F�zEE̵j�z&����y�{�19�[����)U_��?���	� �w^_�"Z�������I��(�G%#����Ĵqs^փ��*Ė� �v�K�v� |S:jef*5j(�L��}�ب��`�`���[���[�sn���m������7�p���X�Pts������AX۟ ��&Wh�������a�`���������G-��$ ��ݿ����?�k���y��������c�m]���I��Uh:�7�k�Ly��bo�VK�o���`|���`����+�
v��}�%��ᝎ띋�6���`*�󔋡/!{��J��U&�b�+�cD��[���T5+�����£�W E�L����'"���!��[�m>����5�v8�����i�d�vH���Q=Yj/��rYҞY9[��P{8˼���Z�|�7nsWe].�1��E~eć�A&FFkH<�qCaa:��� �Wk�(���h�z�|��Ƞ�ȑ���I+���8b:d��G5{5�U�4���XSW�L��#>�ˍ�R��ߏI�a��N\�Cԗ�^j'�.�{WG�tP?��!��	���EK<�6ח���ӊ�g����O�@h��d�/W��xΠ>G~�h��X�ϩ(����p���3��g_c��-'`���&��c�%+�y� KGm����P�or�P}�M�r���~���"w}�z�ਐ��l��v��ՇO��e��d���8��S�ܶ�_X**���DH�,��i'3@�����>���x:�F�
X�Mj��K�KK��������ѫ[��̢��6��S�x�O�/�]�em��,�"��#E�4R[�%�E47Nc�>�|XKZ�����Bi(v݌|^)�柽�#_{���X얮��57�U�14�<��*�i�rHn��"o�'a��JÑ�*��ޖ&���e�5r�rF宲�K~Vx�ƚ��q��%i����+��E�P�H4���uިQ鰔�7���-�s�5^�@8�gk�p�/���|S��s�qx���V�
(����r=�GF;��mYKH&A|��)�I/�BP�0���?�qS##H,P{#qΓ;�@��r�تO�y��k�:�]Z���9��>z�%$�fߑ��41�V�Ut����CV�78�n�6��ޢ�S�8q�t� �D�]u�;�Hb���'��οՍ�9��7�b��_R�W�
��v��Ͷsd�">.���+��@.�1��_:z����p��iQ|�f�?OmǇt�(i�9�퓬�N̙�u�j��и���duG�\���6u��g�I���O�[�����ǣ����\���Vɦ�ϱg'�[h�O�j(��yx>L&�F�cZ��S��h*-���sOX$���͐����n݈���m����b?.�EW��ٶL7�a����'M(����k��e..�?�EAK��0N�'uoV���v����Q,�&�M�A�uQ�_�XE����NK�hq�X���mh�d��fxNk]`�0�D���g�P	��OxU��ˑ'�5{�&���n"����z��5>[O�Z�����d��]]���^���Z1+��\�
�����J9��'\��*F賄C���iJ�G���cƭ�W�+y7��Rl`M̙���;������8��Ì2���!��I;��U+�}G)~��@���tU������|�yRt���}����:DJ�kY�v����`��y�b�4ݠ�Kџ,�c��}? E���ѥ$|�mx�Kc0��e����̚�E��)�tH�m\>��T��bh���ǭx��W��m��Z��:��h���r4�7N_����h�Ȕ���P�|[��OmQNȨ�y_�j���U3:��
M����q�/����L㖻c� ��Ju��v�sg�����i�������A���	��閖�n�f`��y���}O�������u����+!m�
ȇ�"E%�ScRz�xZ"��)�['���tߙ3��.�*<Dʱ,/j���9OT�I)�-�X��[��u<�@�7���<��Jh�m�� �`�Wwcx{r��e�K��j�	Y��Z��`���</+��L ����J�zvq&�4k
���԰��,e�9��n���}��+d�`B,h?i����zL��y��}.��Y?����ZND������
yJG�����V?��)����@%�+ZHx���c�E!m^��[��{�E�o�/�V�c��lI>�_a*�Jx��?�򠺢c�ǧgy�.�,7��y�ؠ����myCnq��f��Ő�.jb�K�Al�yՏ��Ih��l˸S�]��3��j[���m�R�zJ�7�^�myQ�q��4��P������?8�.bP��!8?��b2�\ٿ�<d E����9j[�|!�vr��Y�1/�43J�q�]�6��ݤc�&�6�����JLgEj��d�i��(��j��k@~x��ㄮ�a��l�Z,�!J���� 
##}r�$r[������ޮ�#!��C��}�f�\;}� �����e��J)k[�rԐ%O��0���NCo�/L��<6��a׃�VWf�M�%��s}~.NfH� B_ �ٱ����1#��e���S����.���%/��I��P�Q��'���r��n����m��x��|o��1z�1'}c�L@0.!\�������A�,�,�4S��or�cF�2a�:�Z�J�`���-����NƎ�EE�P��3d{���H8A����� x��5�}bz�����<u�?%����Ɋ���c��X���x���z���:U�Hqx4��qdm�<��Zs\��
>�6?	H�)Z���^=
�::w�S���&Z|��M����T�R���~�H�}p��pyW�mc�~'�^ߖ��mwAz
���9�[>,J���*�+�P���b���\�187�2y8��V&a���ZH�J���vgn���bӸ�a����2��N�!��b������!�<�/g��0���L��o��� \��SK�oLگ�����o
f�vV��:��#t�,�]�9TK��Ur#�%:2{\0����y��P��J������d{X���\y�8����f��T<hB�Ȼ��ϓ
Ç*Ƶ����G����BYuRr0�w��h�sY˨4)�����wB&Sipl��g�u�WB������/��[,�f8e���1qf�[Ɖߡ~h
�c��ﲛ��Sij�g���,�}|�ܮ����~朶Z����װ%�/�Ur��mG-h�ڗyWf��
�gg�ɶ�VA�Ŗ__�o]����c�O b�:�_�a&c�@��Wi���������^���K&���ӔԦM���{=i�tzs]��=�	�f��uMQ@Ec��B-d˶j�R��)2l�8�y�y�[���e����뺐��[�ѓ=�����gf��[��Mvm���Il ��}�=*�°L}|}K�߲>�5�J��;�411*��/C��B���kj�ң1� �)o�!�k+\LײB��������t��R>p���񇓧$��ޟ<c���<Ձ�,p)�<
ˌ��5�.�9��zOUQV��I�"f��ybC�$�t9g���i�&�0�c�ɩ�}��vmM�޼�*�Z4���2-&��e��d����&�u:8�|�b�b����#?̎6����cZ]����U�X�[������x>�]��������ĮaI�Uo�0�9�,�}c�)�àKǧ����{;e�EB�ޡ}�X�h$�����bs{��u���R����O�:j^ w�[`�k�x9�%�����4��ѹ{�Gt�wFc�&-�h<��:D\�H���6�;�i�"�9;�᫯�!WG�/����e��N�����'-��m3���(�����?�5�noP�R�P}�)�zp����}���>M��&��Z:���i��b)D1���D�/�vVy��2!4i�
[��q���h7�X��!�yR4���nfW�>e}|�+��KSkeūm�d��HPߒ�$)����7M~�guE�-c�cf�ѯ<�!�Og��VtF�����+�	�0�k'*x��$�����p������M� �������V���5$�]�䰼��������\�m^Q6��:;�юM��k)|3���̆h�P]�gt���A�I���2/���-��<L׈�����X������]s�A����	J.R+�௟�r=�+Rd_G+~e�/]b����e� ��kl�
Wc�\5}���M��������c�R~�\��ODPF~��o�/6�����8p2��(�Fh<[��\�p���F.�l��rN�d�k�N��;�d�Rz�-��֭���`��5H���+mʄ'֬���e�'���Y�^��@�yU��
���t�-9kyCc��|�
�N���)���5dh���J:��O�ڪ�w�0�����h�ԁ��esrup~����S�ܽ��ҙ��{��y��Eݽ�J*���ʝح9	��gq��ٞ��	h���=X���2��4��؆NCXD,c^�Tq�>�v�E��#�4���ux�9y�KO؁���򇝟��5vm� գ$�6ֳd��Ó���$�S�����Mg�4���D!S��w��&WY��-��Jt��<���'^��*A.r|�w�q[��\���Q&�-��𲹿�o�B��1��W5��Sa��2>�VZ�b�t�b�n����A�	��f�<ynHY�i'a�x���:���r�;�I{��#P̫�f�n*BYA��6���?�\�@=�����.������'&"L��,!��5�T�����j�Wq�����㽪:D�t:�I����D�ۆ�� �C�Y��������ӯ<,Ĳ�/�tdY�������\:�0>����E��@+��%�d��3:%x
s���h ��>�L߼���ԍZ@�>�,���S�і�B4��:�Ւ�� '�I��c͸�&j�/���G��c^טʻ���>�ԁb�.;����꟎�_9�q_�ⰪOdaQL֟V���A�H���q4��v�g!h� �k����>F�̑�r\�<۟�[��X@*"ך�&�T�є�)ש���Q<�PM�5�j����$���ā�����%y�|bCQ5T�p˵x�Rp��z~��-��
�<����RP/�!�o�<p��_Ɠ���K5��3�ۈ���Bܠ��O�%��Ĥ�w��!V���FN�v!D���:�~(b�����$>�;/"��.ZX|���@��c7����dO�mI  ��Q[@���; 񟅃��w�l6{�tm��v^��oܴkU
j���?���3��#�:�`��"H�}��7�&���G����o�qM|�E+�%,�3��!ϓ?f.���W���V���]'��E�$5D�m����z\�:�ξ��{�ܷ�Y�w٬i��|w߷h�÷.G'���b���3�9z�g��0�5TNƓ���g;�t�шu���ߖ7q��F,��vOl^��D�f��7�h��vJm�@�����bڄ�w�м�L�Tg�-Ugs1z��R��6�L3֖����UE?﷣G������9��Llŉ�P���9u�Q���F��P��|�SȽ���-���g����ﭷ�H�髓j�Wo�JG�[�<%���݀�9��b� §E�]m�oGⷨ&W~>��N{������܈8�>I�X���*�����Z�B���	��n����A�
��_�������{?���	�ҽ��y����_$������,�3��sH��tѓ��%�s����tf}�Ɣ����n.h���ǩ�@Ky�	��dx�#��P\qϙ�Xh�^'<�=��9��Jק�Y!���&�P�˂u�'ו� 6�Pe�̏1r&pUW�n<����M���� �����NN�wO�\K����L����/QQq�֘<���eu�����1^�}�?uh�IOt8�˹�R�r�a4��Y���Z�G��cYD���Kd���x�֝��@�d2�u������5y��5Q��q��Q��o��47b�����f��CJ�W�^k�����hDȻMxڥi��3��%��l�B0��x���e��"Ӯ]��uA4ӳsQ�7U�ag����,r����ٚ4�d�=�K�Œ� Wu{�<�7��Xc�J3H�խ��>��2FOu]�O� *|��޶�?���a��۵G�����z��G9b6���
G��@9�ۍ�5#�;O�٫��f9�� D��U����� ͝�*kC�����tX�WPP
h�=g(�`�I�SF5P�[�rf"�0�H�Ru.
�}@�
��$@��.{�mު���p݉��k��+j�.B'd��s�k�������5D,�\M��ɼE��Q��w	>���-���5�H�&�r���"
^?�L�6���)#�ծ���-3�be[T��2� �6��l�l���^����)\�Ay�Ј�x���õ-��:��d���H�c�����=��;�˰�����IiM��K&�>2��|ũ-/ه	s//�v��K�4^!� �Nm�2h~�g�QT�l������!��*���x⌾�Yu�~Y��x�-��U3�%�����?t�p��8jR+"��{���\OSVۊ�f�
��5�:rq�ٹY���utM����%0�\���nM�{d3�����i4M���c�
%x-`e�UJ�w�MC�{8=�C�\�0�mr�[_�U12�U� ��~���!?���!q���qP���^�h'�Ǚ�Pm{�p�tU�[��7gV�����@?(^ t�~ď6�5�y�������e�OA�*b�'8�TA�[����a��x����l��5����������,`ȧ��f��/;y�g�:6���?	L!��`+�c��8e���	�趍�D����_ �"�����"�,[!�1#���}֙�p��>u`���w��\���`b��;g!E�1�8\ۥ�"b���3����y��Cy��n�ڍ�ߙ�G�Xv��Xݙ@{��/�>��Cx�(4�!�L�;��M/��+��L�5��yٵ,�e�������t��AI~r/�Wm� �w&�͢#FyM�4N�|G/ �"��Z���I�FEؿޡ*�*{�����+�.V�4��j
����la�o�|�'�.����w�sUC�W���e�nr�Llce��Q�6楨aL���,:$Z�#�C�!�$ԲA6�
E��Y&���?���R�ܭ������=?-��ڎ�cg�P>$�����B�`/a�pd��)ťHu�-C�}`ֳ���tn��c+�����_����+6�����o�9}CXxt�6���N�;~<�OطewX\"�g(���&a�,E:Z��| �~�B����ηΈ����BƷ�B���anD����Z�?
�0t�[��[��\L-/�E��W�le�ѓ߉�_V䡖���~�&S�b�)�T��	�6i�MZcu��v	�g0��B�xS_."�:��X�k�����\6x;A5>�B�Ȯ�zXo����\�R�C�^=r��}Û�aR�?6��j.���Uː�;i���+������"��~5}�@g6�gy��\��R�3{t��G�2�e�R^���'�u�~WH�<�$F�$��(�r�"��p^= Z��K��J؝���z��Sj��G)���*�f�W����~_���cF�W�1Od��ŝ�[�j�3���v
+J��P�������*�%�"�L~O	���8�ٟ�伽XBM��&�~�v�s�3�B-=�G-rǱK��W|����'�{��u��ۅ�]?��a��2�5G?ߤ�����C�e���-�"�a�+YYq���i�d_��M1���"	/	��I�Z��4������B3S����"T��%�����<�����V+�����Qq	e}]�Px��P�9�_�b0�AH����Vn���_�I����<ts��)$�	U�48��!����k��C��ax��F�!��E�")�6_ s�q�y�
��Tv3����3=nR��س�䓦-o;Vܳ�0Ъ<�s�w_ݭ{ǮNj�'o�]���
���%�G����=�_3,tⓐ���P�6����h�b8��M���(H@��.m�36�����n��7G,��V
����X�o^��kZK�Uͳ:�3ҩ����0侓s^�Zb/�M@:�a3O(Ec�J���O�}z��yN~Zb�LKL�������y� Ѡ���ʶ�Z�SOR���*F|�Ġ��F�F�`�����۹��f5�������GQ%�;e?N.�wo	C�br�q4�%X�h%~+��5NYG���rcaq>��i��KL�h��KH�ea�\:'ڨ=q�ER�Rj|uȕ�3#%�M4��^�l���Pr�Bm9�l�ۅ*�F�H�2)��/��u:�Q�n"98O:�/l�y���i����}��7�c���o�􄛡�۳������W�Ο��H��o�G�n�[����Z�g[��Lͦ�W[c�j�|���A��:mmmsEvv-^�se�t:o���]���[�X\�ǻ���B�QlM��	�P<D�'x���-��x*�Ywllݳ�U/�ƞA��Ly�t��Zoe�)�O\̈́qv�0�S�4��v��y�Nk)���O�GE�'��H�PJqg�gN���$I;[0�(��|��*��]c�4��5q������&�}�ّv�U��+���I3�(e�;�^����v�:��PJ�������Jɨ��'؉c��N���<�8a&,!|�NGٌ�3��rB�>�ƻ��ح�c��rp�r��O@ !����Si�}�No�����O{��TcG���:5�j�3���p�L�_�c��q���tm��t� �����*VY^��r�m��7�(U�^���j~�R,���$���1@{��&!�7O�"���ü���6�ą"h�P)J^k�ŝ:9&o��ܢ2�'W�S1E�ó�"�N�4$�l��wE�i�E�3T;4x�������Y�=c�x|�PJ**��te}v�&��z�����5�~.�XpeD-��D��<s��m�9gd>��0��Z��2i�ſ��>p��-����ߙ�����s��W����}vĜަ�*�ͽJ��!Mj�ە���q��dOn��#���1M��>Y�Бa��}�e�E��J*K4H�I��?;}���	�eo�cB�E��6].G�nkO'�R����_ ��:K'�jʧ�r�z�pğV�xV����]o*�P��	��+�h:K��m?��,�,��۳�'�d��m�6WU kA�g��(�&@�枻�/�bC��mA�͔�f]��/���%֧�Y	�+��5ߵ�����E֞�}�z���r�ɲ��ف�M���:��F�HT�U�����|�-���z�����t&X�_c9���)��J�ņ�VO�7� 4����vԓ����,ƚ���<s*�h�Y�.�)q��ޥ�(��kԌ�|�˦h��l[������v@���Bx��.���j�5�^��YgR��6I;^��Mv(���]&�����W(B�b��[�g.��D�7�r�3_�*W�eQH
zS-�<�-��ON���&�?�A��	�
�m���(ʣ�;��}��ӽiF>�Rb�:�r6u/��$2+H���@�/D&�,n(]�ڊl��J�-l�Z]�63�����Z�g�.Z }gL��;�>�`�݋���ņ1������0���~k��Y���(�!Fa0�35!5��l��R򌗁�]�eF���*$b�kv� 'Ȱ���.�W�{�/���C"�b�q|�;���Jh��%�%�����f��PR-#�V�G�?r�g��I��֬�f�B3��*��ds�]���u���7�S`�W C��:2�Hz����s�W�o`Q����fR��~]f�k�j���Y����;cQ�&�\������k����T`�Q�]�J���io���]���T�q�p�<MXty�Ъ���7]=�J+Ciz��v|�<��xYv�v	E�dd�`\kϚ��vC2���q^�X51a�vf�*���U����D&�D>�]J���n����cJ��b. `�X5��TG��Y@#�~�ܫ#�#jD�N�Ҍ��YyQ�m>��tŭ�9lA/WR��xMk`&�i��X�n3������p�U-̦Ѹn�m�qd8նg~����,D �E4҅Б�nyz���w6":ԓN�?z�zG��FĦO'��i��Mpӽ�X0��#��Xh��mf~�����'%:y4R���_�U=�u� �!���.[jg�!*��͕�����䃐�_@�@3��5?PvAD�5(l�����4mj��a���g)eI+x�<{!$��ZF~Wg�=I��dV�P�;K���%�y:��8��
��۝��v�2˥T�5�_m���
�zm�����ז��`�d[�f��e�a5�p�TV��4��Ok���Ĳ
�Mlq�$�����j٢�A�`�>���2"�"�����N��β�t���}�] �T�3CדIs����m}ᡣ�#<+�NIi�I:K�8#�<S%�Oz����.I�dȇ}֡GyvY��]D2f d��F��τ7{���G��N��Εj�Q�L?AG_ ^���ЏPX��K_kii����~i3�e%����gGϵ�Yg���_Ͱ?!n�S��v��A�jA�&A!�y��Z�����
W`�Y�y�d�ߡɛ�d�_hW���} zj"t^Jy<��y箿3��޹�K�o��7�sv<�ZKBCcA౷�@_���l@���$^O���6XEnX�vy�	�d0��j�]�-�#���Ԕ�㫫ˬ��릧��Ł#)�H3���D����=|d�ȼ���#bb{�G*�v��A%�6[;e���!�bń�"X��}��~n�j{ ���/�IM�OMs�\]Ζ��)�.�a����9x捳I	5�@4^�`]��[G:�����U��kF�S$:XYx˸(ʈZ�0�"�J��㊇f��Y3Vs��Z��i�_�������̌��$d�H&��.j��ib���j�Y���O9疼��}g�C�֓���f�,�[ݫ�N�s䡼��_��5�g����J�B�C+p��1k���
�� �0V�o�.��Y[���ՌWo�O���ӝ��k���Ws���(�PA�xh�k�V�Т��A��"��o:C>�t�a̒�̼�
[j�8��U�=V��_��(�Z�1�:�P��3��.��m-3���9��>���Ubp+���;>%7>��r�b0��o���ד��-p7��T�i��o����<�m9���h-د��c������9Q��ލ.:,Q�l��!�M�E�!���ئ�B���c� ��Nی�N���(�md|s�:(L˂�=ު[%1C��Д{���B��pq�a�@Ćc�!��&�KQ��Y�"����Aѕ]�/�+���7�k9C��7������ki���
������-�v�`��A]tA�FVfCb\��%L�:����Cq�=��WU�+�-��K��}��)<m�̼��KN��
�(�V����,��KA���glD��'�R�a�U~�m�̬�g1�"��G��XIO�� ��X�ڸD5	���#�ȏ0X��d���7u�\On,mü��m��BVЬ��P�i'$�l~A�?u� ����҅�ܶҗ(�0�.��"�x���	]P�r�y1~�@�� �g���s;�vj�t��9�;b$��򸫵���oF�w�w�K��}Pp���v��
�|�|�5cy�Oŗͱ��.��r3�l�P0������t�U�� k�"���Y�&	�G Z��;�C�e\�%A�"8�sjꄢ��C�_ 18�˚4�v����E�<Ҳb2�Ρcf,A|tH���4��І�i����d��B��M������F)�~�5��X����X\���KI�Y��:���^����%kFo�u��*���>�zW5;p`�n͒Go���Ԭ<��ո�sy��̫�W��������V�D�K4��?x��L�;V�"�V��aYUc\��j��R�.�'�Eiѻ��C�N24�-ɮ������_ �qu��;E�YXȠ�Sð���ϯ�/	� ��5� 6L��3��*j�@�}�2�m�G��\̿��o�d��π����l��&Ƣ){U���-���k��\I�qt���߲;fg�`�|!*6G�p�s�s�U�04o��s=�D�ԏOȰ�~�k��uԋ��S�հ���9��1X1:6�-����Ж*R�tF6l�"Z��`�OPT�O�v�.���#(A� ���E&�+70]�{�έ�V$��SD����Kc�O[�e���鰴��h���d��x�"�ܤ[P
Xe�W"�3h�h�Ϣ:�pu��<h~����O�5��CҶh!'�$̻V�X�nK3<Z��Ն�t���B �@����v�|Єk�g\������ő��J������13�u'{P�Y���]�@���� ��]�:���[��!���g(4�+�Đ#\�*�f��l�j�w	���1TbNfkkWI���kw���-���_�'�M�,�+ʱ�륀�"œ"N@f�Fj^��z�jZ�bl����;9bβ�oZma�X�Ix�k�EM�C�{���g�����8���	l�+�Y	�ĵC���3G�gZ�A�~\F(�s��j��夥�����$�A�gBN��a������ð�3�ޅ�m�>3�}l�F� "�kB<���=��V���$��0�݆&�rF�����/�i��hM >�F['N�H���,�S�a�� ~-"�J4��X�7~7��/s�'��D�;�9V91�����}K��5�'X�!��GW��{rq��i���p��wª�м1�_�]��Y����_����0t�t�ԙ{dLD�7<"p�6���nb,��(�2iM��"K�Y�Hʿ�Q�pQ��[��Usx2gm
�B����,���� v97��n�<�}��J�C?�R=k�,^)��t�oݷj���i�@�mw˰�>�QǕڤ�<�[7*�����)H+��by�Ce駒�5H"��N:gi5`�^b�9��*�&s����ʒ@�����(�c����[����J#��0U���#nɫ�>�}���{>�i{l����x�K�R-:x:!�^�>Y�M8U���r'�y�
/�Dwҡw�T-����ߊ���T�$9����V8ާhhI���5?z�gw2<4krCu����SŢX	�qC�?�8��ݴ'��=+P؊�|���]jɭq��߬��T�����K�h���Rc�Q�F����|����o1�B~Z���g����.��x����^?���5茯�7�]���Gƒ������ɑIv	4�J����x,yF|��c	�bW���/���5�/�	C��VR�.�;�Z"�v;���]��Y��Ֆ��\'WzN�+e��P�#��cl|�-)ḯ�e7�O3Ѿ���U܊	n�t]帣<<��7ȐM+�t�Lib@x�H F�Oq��I��T�D|J��^Tx��\YX�O�Zf�k|6�k_}f'fZ*��Q�qt�g8��<�x��h��܎�#�.�'lA\��z�^z�O͒6(>��M��Iu�2�L�ǜE����^ K�p��Km������?�^a*��>(�0��+��ᝥ���>�W���C<4J,A-��QE7D�?�x,8G���7��)�\^�yRq��En�DJ��hb�KZ`��1 ��U�e4i)��	�<?O��W|{!�)-��y��=<��.Mg <����J����+Q]iq����T��|���r:��M�G/ <Io��s�R�2�V
U�5���?�,>kp���R����l�6�������a%�v]�y�\M�˗��zZc䌬���P�M�B�[p��v8U6�Xn�^[�A�C���N��e߿2�	��P�'�l!��n�F�rM��1�;��'���G�犗�gE�)���&������!0Ma�,��`g�j������`�����}qW�\0��u.�u��5z�lM��7���k�����/��S��1�lؙ�*�0VU4�ӗ�~]��;\�<Y�:#����*��EK��jC��x�f5ڟ��/�!�zmBFn{�8��X�*2r��2��e'T�K�1��Ӯ�D��0xt�2����v��D�,%LvZ�D!sw�Eſ�^î�5�U��#Y��9�&���r?\����_+��@���Y(b����*촇�_]͎N�{Z3;S T��mT�L�}C�{�.T�o&��<�_Z��v�4�[����=�[���C���n�vq��݋�w.�m{�m�l���`l�CE�2��,�`�n�k�?�z^kw�Րڬ@?+Ѕ��~�W��x���U�<-�¼���;�r�\4s8�x��;v&5S	���\X��놴SJhI)�o�����O��B����60���Z���){_�LtfTa���V��4�-'�+��j+����W ��V�����D�j$��G�W-u�ˈ\W�f*���@�F�Y���
!�O��y�13��_��`��Kէ�q�������= ��jO��u���㘬t1r��Pa"Vh��7B�E5砋s�M��v��"��B��RJ`�Q&��{�46�`�Ti"��7���*�����|(�D3`}�2*vѱ�@E��+���HY�;р��
B�J9s�貵�Rw\��������q6��Z�嶁��a�n<��eڟ^���Uu��w&~�^�$�
����/�nK)ܫ6Z����5�Ғ����9��m�\q>��ehF8���|b��e���M��6�	=ƙo���Y#"��m��xr�1�f�	)RPS23P���ׄ�3��Òn��?��jT��y�mSVۮ�]G��O#:Y�䘡�G·�IȢ|6T��~x��{��Ty0�Y���X7X�Q�"�L�~�$�on.X �\��ؙE�:�YK2��S��u�T������jP���;��&�ST
�������4�$�C�2Vz�͸�z=כ�C��%��n���uy�������Q�F����-�ZvT�q渃�Q�h�'�r5kXU��P���:���%!���h���l�<Z�D�Z�FN��b�z�dzq��#8!��or�S���d3<-�������d���l�J�� XM����
���z	��Q�.2��*(OJ�&�S�(�������{l��Vb�WmQ'� ��b�HVp�8G� ��&/�w���~գӹ��*
�$G�6�6S�'�A�[9�y=)gߵY��}�S��
_7쪎le�LՁ��LaE�4-#WU(��(T�[���g�:躮	�ט�A`7�=vs�[|�4��Bmv�}BF�7,�f����΃����r|x�o��*)��Q��ΛK�Ka���?gJT�*���+o1#�.y��
������.HM'	,�r��_�Z6����V&=�������Iҟ��j@߱���#<㊳�g���En��Ԕ.���|�oCE�q�fW�5
-�1�qEI=7��.8�dX�G,�{����3�����u���2�ɯ{3}T��6]��>�K��h��'�6�g3 �)$D,V�mr��5�\FD�G;�����s�C(�y<=��r�Ԉ>�U��0��P�h�D�����8�;�O�7�P��q���<��l;;�>0+֥ϰ�~�$��ƥ'��F��o�zV7�O@j_ �g���5g�J�~x�
���;=�y-ugڼA�=ڕ�E��:��U���VP�y���3������[#�1���mW��ryCi,vs:�ϸ.7��u?��$���f^㇊�t��ډ� <Y�n��XA�T�yDOMi�2������4��r��V���{�~}K�r�~��K[����θ�#Vyh�4�.Wg��HEC��qS�.��
��VҎ�WI7�2K�/�3NXM��-S��e}�j@��H]�~%��u<����a��y!����\�!6n���9�6����,%�{��l���l$�S��MW~񲲥i�����J�^����\�^U_�L�� �S�YJ�������h�o5RR8!��iV��@]ɒ�ڒp��Fj�$i�1�/ZU��������R֞�����>�9]�<�����͝?��/���'������vt:�i�<܇�R4M�Κ�V����Ɩ����� ��
���̡�S���ዪ�⥑�Pß�StZmr��X_��,�Ku�j���Nc0�R�W�>=gP�_�mP̩e����^kPmӂ� zcq�	S'�o2�J���&ph�`x�O��JmT�X�; �ÚB�-�F��VyS�8�$q�`s>UL����z���0�C:?+����pDP��tg��]��]��g�S[��r�����@��&B�m���&��-;{V6��Eܠ�����q�`8^ctA��R� ��U���{���?}�oE�����^b�2��.j���cv�����Z������p��`5Sl	��Y
-O���6��}��{BrZ�D��J*�q��CM��R0�-2�q-�� n���ڕ��$�@^y���F�l���~�>Wz�V�W(�}��J+��6�t�"��p�~,�ف3��[f'�����mj�\��shq�~/^]@7�h�b�A1����Q�$B1�R�� ����R����-�W<�z����}W��9Q��T�Ir�Yȸ�l��-�k&6Q|� ���ę���](+����f�XE�U����w�.�C
w�ʩ�Rf7A&F4�E���L0���ۋ�4�&�K]K_��b���:z��s���"����۳5�a��jO-�PtY)r
�/ꓭdR,zo�j���5�%'�J���{�'$��%"\�%��9�	�F�5ӎ�lƴ���u�Gй�HQ��%�k�ʗ��g$���2H%�e�$�i�φ�ۺ���%nS�ױ���L;�g �n���	��⸊��bl'!nJ���4v��?�2]MpʏuJ��h-g��~���)�S��x��@�o���D'������dvh]TFčI����̗8�+���p�ލCLR�����@aV�,ݯy��J�9T�lJ���Wq�H��<�v�U�����G�rhD�
��;����~��t2�Y�k;�����܌���Y`��o*�"�AA>�B�].�G;�A�b�����d�0�ɷb>��#\n����U��=��7n�N�V~f18�no�w٥�|ʔ�a7�d���7�;�v����?�q��*D�HH��h3�>��?�9�r�?�Wu]�+-N鏬�p�f��/�
��K��[��B�ײrcFG�*.(Sp���,/eSf����A�1\�\��߰�e[>|b����.Ќ�y3�!����δ��	pq(��/0�ce��
�/)�S���Ny�rjˏsۗpI�� �s�z7��#-|�/� �hF��%#�-0�mn"�C�a����'YDM��,�t�gB�HiK� �L��r�)�ǩ�)>:�eyҦ����v�E���_�u�?�v\?����N�,��;��ɐ��N��O� hE#�� �
��+N�������{�i~+>H��W0��M�v<|6i��y�\/�礚��%2D1�J	�.ν����G�Z��_̑�h�*�����M����f�S��ݪ��5iD_U��OwM��ǹT����:�j&���6�ec ����_��Di�RPrkJ��,�3�,W���5����Y»��[O��xw�s���Jߎ�eY���b�^4éc�)9��B]�
��ݬ"�z�n��R/l<�m8��y�o��>D��?���͞�d��Ǫ �D�.�lr%��ԃ������S�wS�y^$&�mBr`�8�[�c���N8�m�}� ��w�z9��a�]���y��<���@�LY&��yЯ������C�Brž��V��xJ�n�:��v��#�I6&��_�S���
Q�qX���{��Y>��{�沛{�2�a����/����g�uٰyn0����yY�C�v�3	^;�d��%A�)��HW��v�"D��Ey�0�,�z\pV�
���2y�O���Op��ϯ��@��5G���7��
+���&��)���nt�T������Yu��E�:-���K��)ŋ����Np���{qw����,HqwAN���'�sn���c�=�z�c�,�+���у��<���?��5��t�t\�3r��â0�O�@%ki��_���s-���#�a:ZS��"=�cp���r��&��Dh	�w�`0��*�ة2�z�i�,�y��=V�%eH{�����Ʉ�i�R�`�bv�-!�y���Hd<�uF�}mR�|���E�M����I�+ �
ꦞ��d�Ъ��S"��2,ߧyI�1Yef��3�D��"�kѣ��3��:�'ן�R�9l��C��� �¤6b儬v
���Zuj{�?p,Rwb������;�(���$���qV�[��u������}�9)F9��N�ZwF�Ɛ}>:fm8[Sm]�d"TuygD�th�����]�d�=㱬�sq�R��溪oU6�(����i���u��}�B,��j���:%��Q��P���� 8q���b�������P_	0�)q����ֲ�)��N�D�Pɮv��s�^�qiw�ſ����νs��K�2�;ER���vj��	�������4����ϹA�Fv�S?A��H���b�5��.a%@B�7�Fm�}�����}�*pt��Q�;o������SH�]�#����kƨ�ē��� ġ�����|�F�Y�	u��^os�r�X]�Jl,M�������1ǂ���5���I��B��6��L�OE��R�l%��#��x��l�y|:|fT?13f�=}Z�^y�O+\U�|�7g�r�o��a���l����j͆��<ô͊0~ŕok!���⪪G,���yw��nؼ��g���J,#�稏fx�
!2�Pt��/�����
rΎʄ�5՚���˯dI���^~m~�W��,��	�N892��VeWG��Js5���Cݭ��|�U�S�g��
��[��-������e�3�<Q�%�Ua(�cR3Y9��� .�e�$�X���ԔĲ��D\�:�-t�N�`���K�Ci���|ڼT�+���}ݽ�J���_i�(/H�nS��2���}��K���P�_ZNN�<��W�� �钊6�Wie�qU�Hv�Z���<�� �c��(l��'�d��!�:�*n�h�m*S�'�ݻ������tL�[eXɺ� ~#��:*���5]Fo���5S/�����ux)�<,��Uw�� ��_ ��gE�
����ޛ������ j���Y�;�d)v.�����@[ԋm�.IOH��ӫ��iRV- �4���XL� Y�����s-Wr��IrՇ^ z>Xwҏ�%5�d^r5S�/ ��I�Դ^�A��1QBQSv�$K'£�d*��ģB�Au<�s�#ﵶ��+��w�<'*Y�A�
��g�E{V�o�V"�vk�����3�X�c���{��9q�u�\����0
/-
y��\����V�)������'J��;���p8�:k�h2��U���po��˓��x��H�q#U�"?���%��ē��q_�h�m=�y���;�],2����ה�D��q��$�L(k+-���d)���;���~qQEE%�N�e�-��yꔖ�Cj�C�mEi���ȳm����DM+�o��wG+�=�vt���1��k�j������n��9,=����'��T�o���k:+�iM�I�_�^ !�7���V��iO*"T��@����kX��Z|s�l�������-;mtqffwF�W��V�rd��S~��j黭��++yT$�a}ן��B�o�~	�[��f�� GF.-^-���/���XL�ŀ=o|��q1le���}���%��YO�5��" �����U���8M�y�5l	C�{}�d�Ű��#�p0�
���g�nU��x:ƻ�B�/��A0��SЖ;?�E��Dl� ɀp���\;^�ME�7����C��¹-	zdJJ�^C�$$��,���>6�o���{�RV�D���e{rUPx�=�;��Z�A=q�ØBx������>U��������9)�]'ʙ��SZt���8���������"���g�u��gA�&�f0�C���j���R$\�C;]M�
���P���,c{����x3VW�5(��睝?9hl��B�f�r왙7/��7�Q�]�y;��[���Gm���B);w\Yr��&�-�I2�%Κ�2���l�U�t�ڙ�N�ӝ�	�����|4E١ܧ��`�˂�`�_?^�(��rp ��^ 8J�^�J%�Vr����m��n
O�ͳ)���W昜n�SK���!(/)Ebz��5�0|0�ʮ,�b�2A��<$}��:)	�&��c^pC<�AU}0�So\T3/���BQ�\z�:|�/���B�Œ�=����o\�,�1Ǎ~|p�E�"���z���X0��E|^�{z�%�it2��� f�������]?@NZW��Rs�G�iT�h��X�������(#t��JEB�����)Y��u�aƃ�*�(S��A����Bh?�r�j/���<����{��t�e�I^������}�-��1��$EfE�=u�8�8 ��jq��)�Mf�� ���)�n<�9�5{�z8T����ݦ1�Zo��֐�k����U��	��k���� EN�]3ܿv#+{���d�Պ�f��q�6����9�N:6�|�N�:K���m\�����i���YDϳ�3��jʖ�G��^ ��w�!t,$��[k���&O��c�aș�-9z�5���Q��?�ڶ����,�Vy�c>�}�CO�[���\��ǩ�' .���mE�!ټ7��c���L�?��D_�����N�<�y�}�v��M<�̑��{���'q�!���;��;C�RӅs�@;��~i����b$MO�<D�|~'��V�^"�|��c���S��3���r�߅�\QF��I{�����_+��)\�"��|�y� n
.l�Sp�߮V�'~�����/�9R�|!Kb�(���t v-�(�%j�B4���Y)<�X�N�<���vrB������ ����`��%Q
������n����&�Up�WV]�3�ZT���]ğ��U4Z��Se"J+,�5'�S��uU��0P�����F�=��Rox�+,*l�ojvu��GHR�@O�5z�+n��(�/I]lѻ,����Z,�xb��9����[x�����8���;������ex������)ɞ�,�}%�4��|�}o^ �'9�߹I�]�V`���Uu��hD���U_�~F�D�,au)$7��>S��]|�����h]O�`�L�.�R��2�e�q�S�U��s(�\
؆�3ʶ6Qk�T��-�=+�"�a�PPW)����'6���ɖ��|B��U�2��8�O=_)��dX%h�H	'B'f��U����2pW���>��5x�|�D|;^M�]�.�	��Em(�I��}���¤�.�\Q�.}J��{�`�m��E,����4,3� y�3S*86�C|Z!�B@�<(G�N�A'i#�!p\�.#�p�l|u�FXAE�G�o?&K��HZ|�	���y��S�>�͸��Jx/ v��5���"x_�i�ᮛ�lm�v�J��m���6�-Hc9�v�4R�Hd����f�w���w�%�	1*8�)7���^�ೲ^
��".�,"6o��ouݫ�)L��^��s�m�%�0!����C��;�婿t��+��j*�[��V���X��i���^u�c]�bMO,

�b�A��S(�����<�5_ �z8��]�X%,_W��=��qp�4�L�̿�lŲ/ʉ­�̝�M"���~�j�Nɿ�8�&�bO2UyS"�h��m߲K 2�~ V�ʷu�N�h�11m��ő|��sM	�wLD�t�
KlD����?T[���$���)�W��?V�f���їW��ʺ���;��*��;�s��]j���7\�t3���k��8d+�Q͡˂ v�������y��:G�6����^�hH[���������{�?Q�{EI���5��qS�ˑ�15��.4�>�5��7]� ��S�Xp&�]l�TK4H��,>T1�.f�����Q�~Dhl�-I�C��{���f�:���|��ŹKZ:!��׿������ˤ�zg��ȯ����̼��D�[,yf��%���ʂ%7y|�$\SS�]Kx[�ZԱ-<�E'�T���DI��tO���S����?�岙����S� xN'�����<o��G���jJ�VE��I�ò%�'M�2>����ͫl4����uq�G��)�N���j�\
+��ǆ\�6�]�u�����0+�n�A���]u����8[�+�@)��,�7��� 	�ͥTd)��⨃C݀���t-k���ڊ�LJ|��EGH	��u�J�
���[�nN ��f�h��Qu���k�!���4�(���W}c���C���i� �֠��xn�u}ˢmB��������eU�`��0FoK��&T$w�Y�M�\=�Ǵ�֬�3�?����OIw�v��`�衼��bd?5u8�^P�^��Y�6W���4�(���#K����1��?��惧�S����������������]�c.:�y����,�U�U�L�]lø��"�T[��m#���Q�h5�'J+7�Kn�L(�+���d��$׌��!+�"?����\CRA1���wl}�1�N��n�,���=\]�q�prHy�٩K=�dYZ�"��hc ��с�6۪0�(�PN����A��Gߟӓ�'B�("xg$��UeMn�I��w��#`���om'������\w��Q��G�}��w�Pa�K��Xmq�32k�4�9xW��V�W�~�Ċ���T��v�Z�`=D���-G@�K�L[b�&��Tzk����}�(C�I�.ixӇ!���t��hU�����%|`k�r��e���ۿ�����1����E��B���mw�b�R�[D��S ���9~������#�"6�-��NN^_O�y��QSѝW�>���;eB�㴢Ļ��p<�P�5���ј{&�B�K1�8�]c�U����'̄�$U��'j�mu�n�~��� �(#�L=��Z&�VWS��DF�OV҈pZy,?�<c�Ԯd<T
�X��|��VRQ�)��
����U�ƳZ8����mf���ϡ(��Wi-M9���V&��̵1α�F:���6.S�=ZE2�V�Y�Vz F�{7J�϶�=�Z�T�"���(��*Y��j��C@G�/UV缹[���ZR�U�Q�W�����Z~Cp#�ɸ(���|MM)�ղ��C�ۡ4V��c�B���}��qx@�S���?p��q������Y����|{�w�B�����Ü&���T���S���H�Y� I�}��BU�C�о��P�2�E ���7�Lm�}��w�/c_��(cT�#��KX0C5��͠,��;rڿޭ��Ӹ��z���/#_ �Z0u�T�$-�� �Ƭ�V�H)�����U�C]m˼��#���5�a�����h�_�}�d���Sl�8.���YC.Q���Q0�:;yIZ���u���������;�v�bw�#eYS��}$�*�SA�_�J��l0�/��+��1�Y�5�Tݑ8�M�U���7������
�h�B
�����Io�'��D7(!�g���P}!�]��:��r�P�O�KpR3��z�l��h����oZRm�ffg0-�Ą�<s���j&�ն!x߼�� ��3
��h,� �T���#���C߈ƻS����ڈ]Su�R�Ɔ*T=	՝O��jO&�;��`�t��s�?>�Ԑi,�|�2+x�XOq��q�"�HR��I%?�	q�54_4Vqf��a�J=��`�
U*% 8}�x|��-0����茔}qCd7����I��a�X�苐�O���sd0��@T���2� v�G(�I|��Z�&zdA����P���{җz*�526��[�gh&��%TO|�����Ď^ ]v�֭�]N��Mc+�5�x�B��Wc�J�������1_,W�?��vJ���]5�̦��μ�3��,����>ᇥ5֖Pٴ����Y-+�_�P�I�#�Ft��V0 taT����������aK��kkl��bڷ�P��G)�r+K���JS����5>��t���z�[V��&���Z(g�ĭ�;\�PJZ���j��V;ͥ���n���ϴ�f�PJ�dR�P�t�nR�cn���JMW؅��	�
!���5m���M�P���U���&,{�
�|�, ��TXN�ũP�/���S�i(z�������k�|�C���`o|�t7Wa�+:=�`y���>�4�ݿ{[�82�9�����_U{�x�γͯ�(�hx�؟NW����g����t��)���A�^kpXmJ2h]�1�Z���45Y���Tg�lv����wK|�������:Ӷ���0n�Jg��EF��2��K��;kϔ☑�<�[-؁$�<5zM��Ω۱����^��Ҋ���g�����}��I����&*1��Ƀ�6�jtjF�hbe6��z#�Esۃ��fZ��M�ƻ��4M��]������_ 3��T:+�����/�Ģj�JGu�$���<הR|�П�DM�TR��\R��0���w���v����\�v8>���.��<���LT��8���=�氡�r�RV^w/�7TX�N%Ru0j����'�@����J�'��[^{�B�1�%Ȗgƞ���G��ut��ӳF�j3��	(�
޾))�;u$��H�i��OMv��=-����V�nAO��a�|ԅC�ƣ�	����D�
�~�ؖIS�?�A�г�Y�����!����\^V�l�Wf�u��������,E�� 3�M�~|8��pM��ƅ��l/������Llp����gr�)5�>��<��GF�<����G��`�����������2ge���7V�����������i��095�l@.E�&NT6W�D���ޫ���sH��1�V`���<��^=�!
)X�
����A84s��U�~�4�DB[^Y^�5_Ip��1����l_��`�:����[�I�D���-/�"W��q�w��E�k�����qN�x�o]U��_UCeK4��bF'"P���-��7�+�*ܢ���O4Y��zOy��"��a*�叽"�s���[(B|�	g���s��sk�n�uG��k�*�x��o,ᒭ7/��0�4D���Zj�֐�����|�����rϩa�I��n&y��(d��e*���w��5���^�l��sr�ߎ�$)+�����Nv���?�Ynvɰ{�P'���@Q����e�8�R�4	��j�A?����d`�5��w֑��au+���b<�I���v|t��HV\�`��)�S��6��	[��}N�q�^��{S����&�-��~Y(f���	hl��[�jo�����j�j|�ļ�Hv��3ih�R�*���[����Q�+H&�W)I�T���fGYzڣw�f�ŗ��(��N�����ƕx+Pf+�kVTc/iE�!��L��o@��I����͍����<�|��'�Z����4 �2��)���S���:˔�?�(�˰��R�e�$k���2���YnyZ]����7�g�f�g;D�JN����<��yaV��<ed���T����[ـVN<�����k�����4��߻�Ā�
^��p\�`\�/L�@�=�j߻�Vya��v�/��ڤ$�\,Sio���b�lFU��>��R.�o뀴J��wRՈ���RS�r���e����$�
P�uą���,��dO�آH�'8[��˱�1�|(
:h;�(����`����%�_ii�铸�S����$O��5aH\��aɭO���Q�{��Dm���s�:�Q%�$�����;���M$�k�����@ej|Q�����c6;Y?����.ek�TQ$�$|	��d����L�A1���Ab+]���Z/(Zv�0�Z�Z����C4�$i�0��P�j���k��J'�W<$�:֞��.�m��c*�
�* eηaU�2ITi�^��qf>\���{1}�7�Nz3:�k}�p�!R��頱V�5RS{ƂAߚb�ʘPld�؇���W����	wmIvl�)����ŷ��*�v���e�����kp����1�1��GT�B�ܘ�\	�%�h�z��>UT�>���1�.�������'ڛ�س?��W�|ZYZ��7Ke`$����v~�!$ȸnԀ��N3�@yE����r^���_�
����*�wr�v���b�|M3��J;��?o��1������� a���#ֈ�ޗtn�u��q3��f��u�Q�HA�f�kF�r�r�4�=��k�Ȕ9}��_���<6�%�m����e�&���c��5��#��	#�n1[��Ւ�q�����s���'X���+Ү��6� �"'PQ��r�Do��Y肶�Jη>�lL��8�;;��̄TT�хe����%����Y�,�aĵc�����&Pz�neA�k4���������.U^ Y/ ~y�˽]�ɼd�9�2��VOyw��5.���)f�Ȉ&(vl1��������onXi2A�Ɖ�A��/�1M����:'�����2%��l͆Y]�L��~�9��X/wȑ�S}�}��5
ڭ�~#�+���`_�X�*��g�v7f�m�!�,�S�'+=Z����xl��<���6/����v�21P��$�v��[�d�e�[{c�N��1S#��,T�Gu��*�x:/(�w8%4ER�ͯ˅�+��]9������ ��Q���wB��l���#��Ā8}��ky�}�m��T�`��!�g����c�?�$��A�k'��hw;hQ?�69�H���AC~�Ո�U�؈+���^�d99��g��V��$��I|������s��;vL R�������M�D�����}�G���i��Q���q�w�i!���_*��Jc�>n��ٟ �Rw�$-�WS�u9|���}�4}W��	��_�R���e-]�騠
��=�6�8;[+�Tߊ����Q�\������͹9�N�L�]I��>;?�1�ߡ�0	_�X�4����d�>P���;�����7�T�(�?^��L�W�:c*X�dq�uh-<�1��������i)o�F�Uu�o�mQ��O�
�m�����o4��C��+YW�U�K�hx�FY��������O�h>JT�2ɂ6�h�g�:|����!ӗ�w���c;q��	-*]�Q���p�|c!q�NS�xE��i@���7S�ҷ�1��f<�ç��'wnK��MH�AQ�[��gE-�YvĆ1����dd��-�`���z�ir��ZN1C��/ Dn�L�UI�kJM~Z���M���D�z_���߃v^���Z'��x�'��ۡ6Şs�w�6�����^�r=���C�q�F��w�v�(�L!�_��D�y-���P�\e�b� �?�7~��I��iW�}�����J�l�=��P��2�V���O�[�~'./�s�Ք�AN'\�y�bC񢍝XO SoT.��fhD�P�>�,T�ʆ�p�26x��woi��$�)��X:��.ܷrV̶�*����z��W�Q߮,�u����Ҝ�4��|�5�:��N���5���R�U��_������;$̳�˻��W\\O�1��~G�֛胣��-pJ����бsL�z�Z�|�A'c��w��g	?ғ�V|����l]�\����|;�2Un��i��z  hDͧ �E�mr���w�W��R	oXJd���t�L��n�ee��%b,$n��7�Ɗ�ԯ��斎M�*+�N��b�v�bZp������Z�E
�� 1!�K̩�ۖ���fQa`�/���?�iF���}�R�ت�K���͟{cbfS7Qm��ˀJgQ�����3�2��	�50���?�Y`Ĳ������k���^���1F�Ʉ�.�#�g��R�����- _���H�Ed�qA�}UUu���űT0 ����� Q/G�g�a�W�U]�I�����,]���#����+�-���*D{����۾�lJF�t��z���Nb�"͠��I��7�Y9%#�;�&�Ys����Cٷ�����p�4�bM:k m�ۖ_�Si�yv�<��Uv+�m]�����5�� �\V2LP��ݸy;���w�C�C+�V�@޴5rxNY��>^���u�Rr���߼2�z{I��,*������U�FD�B��r|��;�9FJ����g��|�D��{U�����r������V���^hR���(��Oc^�ZA�K�Ii���
�}��QO��3,����������I�P�ԢW��-`oM�=����ZR'�2�+��8��E���?M�	D��<<6A@=.���N����]��7i`I�C�o���F/������l��q�m�� (5z���m�� ����T ��E*�H�6�?�Jɞ���g��ۤ�����g�UJH��Ҫ$W`����fS�fs�Wk�����t�d��+������Xh���z�KxV N�o��x�n*�
�\=Z��}I�i��|Nޙ8V�36:&�8��6
�N_*�J�2�����x~���NΞjV{V^�J� �dY�!�vK�i�3K�r���FM����1$,��|��hx�ES��A���G����R��X}m:.�g���o+��a
~��xN��z��;Ӆ,p�XM3YE��(����:�d0}o*���ilo�o�_K��q;�)�uW�hj��nT��O��o2imT��P��D�!��]���i(;r\�gl{o�h��#J����ҿ������$���؇�s�{�
��þ6��&blL��Ju������*�L��cVMMm)��\N�����|YY��I�ns���>��>W��uN��au{��b/�.�"M�K�֐�eC擋+�Zda(�i�r�n�j2.�dyɰo��[2�t̀�v�^O�O� �f�-?�v�	���$ej���mT�rk���{�_ۘ�Z����`���5_�3��_�������ӢO\��o��'��c&>׊:j4��w���>��q*xg>`�OU����Q	��]�u+�s��[�B��Ƞy��XU��(���Z����)Ŵ_�%��Dd��6~I�̨|Ti����H,�2��~��.���O�a`����
�
՝���0-z0���O/���'�v�n�S�:w��_Q2��S�q�
Eu<�p�hO�I�T|Ԣ��
�.�����;颯��T�I�N-Ň�d�״JA���IB�����^�6�;���N��E�R����`��J�{H�1*���Z.�N�sc��"gˣ���-�:D�5'A��~fur�#���1*4�������9�N����č6�F�>~u;��|f˓=K�QF���9��xԄ4�?�5���=�-/	��4��ܬ��R�*�zg���]��g���J��B���W(������o��V�p����1,���6;F|�+8G> W�Cq�ߙ��l�7�T77W���|#�vp8����ٸ��~� ��Y�&��y�}B
�b�n��-Y���W���Zk�������%�o{{E�g(3��'�����_}�&&����7���'�#�n�œ�R[�iaG��-�<�G{��{���A�J���=���a�W���?tv�M�	*���ǹi봡Y+��q��}��77Uk�A�'TM���;��@J�%�ڟO����a���^�l.p���ă>U��q	v̊u�h�%��O5Ы�W'�I/80�/QWKʁ������w��1)����1M��Hwtͤ���ͮB�cF��zۆ�"�_�}b��Rv�z;o��9�,����Q���*Y����7W����m��TT�]m�Ϛ���N)y���9�A�!J���IZ�}�Q�+�d���t�_/����_���r���c���|EG���_'K��X�i��0L�|[�Ox�'�7M�Zy����`��r�H�h@��~��~��?�޺�ɉ��H�⁇:6�a��ܤ�{[�l��$�����rs�^2�4�Yv��Z�l�
E������7��Zf��h��#4��.��m��U�,o���S�H���iMWXX��n�X<Ы��t��I����FD�a�TƩ�2�}�<ߒ��;)��q���B�5�O+q)��S��#��6�ݣ���X���ۊה!.p���,����Ml�!Đ_Uy30Ov>4$f��7"{��z�K��S>?(	0�{�����JT�Ȥ���*z�N�Qo�Y�rS��:M\I�<N�����,\���{N��e�eE��!��j����D��D����> C}'Z���**�Ժ�H�]@�v�+�Bf[�\�{���ӆO��g��s�Heo�e�Mv��T�E>L7yŧ��%�h�r�;��2����A�)R#;�S���&������a
e��-�Tw�~�Ϲ�;E�+H�8.����M�[�3>V\H�U,�M��\d�k�����K�}���F��!9#;��s�E�X��D9tK����jՏ��5�6ԾB�@2M7]�!�` ��e��N'à��E�+Mk��������G���yq否Yy�v��g���4SZc���aOO���v
'�wh��"K�	Z��7I�#��k�j����v��V���'G��\V�bxX��r�5�X�=s���ۺx,��~��L+��7��F�������j+b+�����jI����ǎ�<a�ol��Gb��o����F��+��J��hj�㊾ݖ��2>�y����.o�ɑ�aQƯ��v��Zy��|nUI8:ɯ`����%���l�`���}�Ɓ�#\x�w�?��I�z�Gb���
��%�|7ml����`�DDvs�G��k`Z���d��L�
���5͈u]�*4��べfȌ݀�2ο�#.�+JG���H�빞�'���7HGM��դ��}Uֺ�D�K0�`�|p��A9��]��U�2���p��� �/M4���[oX��Ӕ�$��1��h+���K���HC�� n:ȋ\8G�6i����ޙ��m˒���[�L;�qF(��'�*�C��~�pp�Pqc�4: �U���+͢,<��İ��̡��\�s{P�[���dy�5B;�0�-Ч,�"ȭ�b#P�Ƶ��
�iz2�-7��,G������_�]>�kh��m����ʇ_y���i7��<�P��s��{�<2�rmT�],v������15�r�]T���'M^ .i<�2S5���Y8>���T[5���� �wO��A�(�Ks��4o�}��)�-sM����*�[C��W��Y��'�د ��
����m޽ <�V��{�M�țZ.�?v`�BZ'���S�hH?L��s+�Z�Ț�j�H�{�x�L��x��4\�-�i�j!�n{" %�5}�82�_��'��Yb�)�P_��4f��� tG�z�0̋RI8�f�A�kO,���Y�M�$Q<�FD�%��%���jW*}8�d-�IC��5G:��;��S����Q!�J��;���H���[ʎ�t��fU����{h��8Z��S�ZNwG��q׭�{`�F-^��`�=��� y���i���:'���E(�����uħd�$�8����Ӭ������4NT/+�9��x� ���)��ArLҢ�������0�h�S�c�oo�@��j�<���^p�Q���E/���u�ie2оP0D��k=���ē��We)I"��u��)<�d�>To�b�f��G�>ۻs��w���{����j�u�Y��x���c�����֖�=�SP���J/�ɖ�+т7�p#ʞ���*��	r���Tv��h)D�����_'�9K-n���ݛ��	�dc?� 焃$��l�s�����xQ)D-�������δ�f�?�1�N��V*V�RDuѐ|cD�I�Q�@��._ h�Ռũ���h�����.��ޕn�.Q6���ɌP��D��y��ǧؠU�A�Qˆ�V�TV%�ٔY���*���K��t�C�}�:�)x�o�-z��%�B�/枥�B8��1k--(kgp��U"p�x��wI���K����(o|�"K���P�DX�eO��H��-~�&�=3�"�};��"c���ή�c᳄��}�鳘tcw4�AU?�?�RХ,3O����R/ײ�����"������|����e������r�������]4?�:�%@#��,��#=6��C�9���2>����r%nctu��J�
��W*�jmS~XV����5�լ�W�o�ͻ�m7ӷmnʒ�����A�{�pq���8�p�Ѕ<�
ƭ��7F�?F�;`Z��1��=�u�ɳ-{�63�?����L��_Ņ9�~��D3_m�X� ��
f �P�ߔ��S��t_�w4uK̒�z猨u�*f5x�׮����NL�*f����Swk��-Kq�-~U�|������f���#�#�/�u�x�{Ҟ<'juU����(��5��ܶ���4z�և��G�\��n��@���������)���)�"���aEv������b�/���\�vy����r�Y궺��D�o�l�e�f�Ew� ����e��[��%Û���cCQ��G��_'�݊�;3���8�?�O�BW�Ț��A�%hDN�TUMh0��`Cm�U��v����y�"��l0��ò�fB0A��ڲV�:�+r@����#��8.k�'	C��TVR�kAV�4�椦J��C���ʶ¦�~~�7��$�3qK�E��shd�7:j]�P�������ږ�G?�>U�Ӟ��ħ���6�}�P�b�����c�����uk�Kͥ���U��h�N0�|��7�ڔ��"��݀*YS��+�$��A��|���?�1n��[��-��������'�x"�Z��Oc�a"�¥nNl}�?b;��m��G5bxǩ�2Z?rXcZ�K'�S�A+�,�HJ3R��/\�!S}ށK���ӿ0w2������d�k+-��{#�t2�t|ka��l�A����e�45 �.X�E����&�"ِ�%�*<���*F��q�S��y)#��[=��U��鬍*r����)��Ȩ�j���
;��q�Ԋ��1� ��,gnw�B5�3�l�5I��Ęn�sK���jH���<��F;h��V�C3���ط_�!�o��z��{�z��qQk��x���"}}�'s�	���˿4"�W&l!�#��[ib)~>����q;��g-I�1}���z�,G ��E��<��Τ��D�}�v^�'UM�)����i9^��^^����w�����܄z:��p��A�.6��>'������N��]�wI	�����);E�xF��2v�n�g\��EY�V�i1�|5�dw��`��x���$Jg�W
�c O��h��_�Wd����|^W���Ǒ� M!i�7P���,<�Q6ZW�]6Ϛ:�(����m�����|�y��H>���'�A�����^��4�9լl�}
>������5��ҁ�fӬ��8V��`�F,
Kw�H�֓4sba0�X�%�1+�r��C������(c!�J4��'W�܏٩���;����1},��9��� ��2�eb���Ok=�I_�b��e�oޣ�ᬔ(X���tQ�
:=[_ ��^�;�W�����~��r�&�,GsPۚ����f�QQ�7�%�4*�����65k��TQQ����^�{���6�d�<%~r��s�g��0G�u�(�8b��C�t�.�xE[�x5V���W��c��^"}|�5��X�`p*U�s@ὔ�,�f�K�ds}cb�\a<�B^�k;���1b���R�<e���j�(��ږT�Z�]{�X��1����G��-F��e��q� ���	B,�������-*	=���ο��-�F��+�ت�(dDEC��=��F�z�����)(��CKsC&�?��ҾS�\�	���U�����F�M�N�?�dl����W���J0nQ��+�<�k ��������\���.������a�BFddwK��K����*��h?��[9Z�~��9�K=���b�E��~�p��K�p����j�w��m���ܽ���5�{S�݌ �����w��Xk6导AN��򎜻i֦�ҳ���v��<�3��X4n���j�iESU9ua<�ٺ*t%eT�bISXbi�+��(wD�q�y�#1B}��%6I��"�9�fC~j��^�����?�}cw�����4h��v�ƶ��6����ƶO�4�m�>��������Z{͋�5s�=k&��������J��1ཨh�-Y�u���Lj�_�=X�'�L?����`������:��g�m�h_��.�|�P\�NBV��,s��|��b�Һj�Y���}����L�n��ቄ���'��C&戉�B�?� ���bW��I�rpL�	�����[���(k��r��pL1b�-����[n�Z.�.U���)YE+�s�����	�����<:�-Rz�fջ�UX��p�0J{�z��?f��+�4O���),3Y����2�]����]ֆ���� ��G�ƃ��MJӐF$����*��n!�.�C����Q�2t���UP;�2H���������J� 9]Jy1]�<����V�v��naK�w������i!�G��
�����w��	�?0w������C%��1�SU\n-�ot9�WU�7.{��Gw:&VW�I@.�����YD�����+<U�H�bZ�X�DZ՛4E��}��^�Ч:��A�%�6Y����9�1��v��=r5䶠M�6�$�ݔ	B�~1Fu��,��y��0���:���t�E:\8[��]ՖwեM<`aUpJ�sHR7��g͛���2J���Q������ŝ}����["���x��!�q�	5�Vo�f^��<�zlnߑ�ǜ
�'�Q�۶lM��d!�Y��|�Y�h�r��/���~ٍ���	�=s'�W(�)���������_�~�/ͩYY�e�����X��C}�W9�Wu��Y�1��ɘ��\x~��Ώ�i�ܑ�����b�kzr _ Gc��,��^0S}�m���Ưd�\��{�����A��n�8ww��I���E��':o�|u4�/fn�Y�e%�)���;i�qw��n�Sb�&1�ϋ����̧b����f�� ������ڕ��vQ��WD�L�/�	�`}W��d���i�UR��ׂ"Hu��;Ƌ�KK1g�/bHKpͽ3�ur�s�F��4�\T�3��֐w��<+cb��ˤ2B��^/�ٻ�u}��
&9�"���CpZO��&O��W�S9U�g
u5�֚�gM�����EE���GH+�L��#&�*1[7d�u�t����j����Ko�,;\bJ�iT��`�U��;�Q�����C-1}h�x ��������&N��ך�v���Aܛ�=ʂ5�g��A�`U"�^�ПlS�Ƭ�����z���M��BI.	�k�h#�ُ�Wϐ;��Y�@f�-��84�^~�_����
A�o>fps�\��Ѐ�_����"+T"�r��������6<����w�sL�����ͯ�op -��Dd�{)�$�X�`N��l
K#�TjB\�/r2/Jc�����1Zm>�Z�`2V�m7)$��=�Z�*o�X��Dj޽��v5�"�|�dnΩO����ӱ��bQ'�Ӽ���X�l �Q2\�b���Pr����9��
c��� �R���&ڒof-M"��oo%�r#~�J�W�t���?i[ؔYV{ ^�.�8�B3�=�n)�}�F�*6UD��$�ȦIh�D��
�9w�jCm%��vww��ҕ+eR1q��Hh���ꃆvD�����l�wm4���@L��i��ӭ�|>z��d43xʊ���W"�����y���_NN%�O(+�?J�szG�h�C���4?|%5�6���{��yT��Z���ˈ���v�n�U��Y�q��a�x��ݣ����t:X�A��X�I(V����WaƦ��-�p��[�͓���˦�ϥ�/���d��L�H�O#o����hTV.PB�`���K�����������&X�
y#B�uv�� k>;�.��L�:��BF�l��.����,	"�)G����Y¢eғ��|�OZzۂn�W�"r��͕��[���x_����ҟ�}�5Δ�(�
��O����� ���SD	4Ƥg�	�P�]LN��U%�-��
�H?Q���WY�@���M�����r�"�U�^
{���65����D��d;�Ĥ�*�V~��]$�'l&���-�iגN�ȥ,y�*)������4x�'+B�L���	-P�q8��dug��h'����6/���.���t�a�T��Yܻ^��A�s��v�tY�h&�ؿ����8��˸$�c��d�	x�T�x.�)��lp+l�ﱌ� �m��3�)vl�i�sƟ���;��X��Ө��j�T�]�R����t�0TdE�N& #��>R$4�kk��K�26�6Q�T���(ȒY������5�b�pYhywP�"�k)6N�A�&���0%�2� �vs6�tC_�*��I���V���c��N��cύd��r���p�@qzx�m&<�1ȧ�2�Rlm�p̖I�خp���f�?�_�F �'�~�ڿ`��Y���?��^�*S�?N��&�`%d���I�c�V��K�������ݖlN5��ɗ����m�Iv�\�3m�0h!W���~.�~� >D%"T��H�l��t���+�����dN�Y�	�9^nL$��ݭ ��	(�k�b��$�?27�0n��µ R�}>������ڣg�%���J�I%���Ĉ�%��T
�z
��E^�M���_%�d0e�su��ϯ�.����R��!>����A���p{SF���w�3��f��-���p��csc�Y�pV~.�0��|��70��B�&�0��[���ًО���)��g��E�����&7�f�dNM���۬��0'���d��	����H���-��S���v�����n����u:�����%M���qE ��^����bQX@k�����w���H�`"�6v��
Q��,��u���BH^e^Մ�����pҸ�y^�~hBD4vLu@������� PA�(kfh��!q�@�z2f�)�Le(|A�K����7���w��6�F� ɻ�@�1���7٨���K-��O$IP�Ҏ��#G¸��.�ח�ebP��[/�S�-1�(r=c#?��θG:B�i-04뮭���bc2Q�b3�P������,C��x!�hN@q�M���c�(ض�v�1�-��g���=�-�?���2p�Q���T���GC�5�u�ky7/N�14(�Y����Y<O�����Z��Fl&2Ya�Q^Xy�X@s�h� m4�֩�A{�b�X���NB�*E�אjAdB~F{9���2V-��rʯ�ٴ�s$�I��+��tkNc �����";'��5{u��k�&�)��i���@�g����:��Z`���G�	��G�b�)�*� ����lBN��{��)ַ�S&%�֣8��l�-��#��\sfvK.ǻ�7�`>;.���E&hd�r{4�;�x�G�ңC��+lٞ>�'@�hnPC3��8�a�7�+�ŀ�5�=%'~�X@�zE�LP��p�ܚ?*����)Y3î�OL
b[�^+�s/l'U����^���.����۴�:C:����W��5ߗ3�CoQ�=�{�����*�(�����tq�
`��������z�[U�e7���s;/���=铓�y���$+�O���p3�O2@���"1�W���N�W���v;����95�O S���9o6�kV��d@���_O�~�|�ImF?���V�@!�D^�HL�?��F�N�3�_`��
�%�_����!c���!�ނ�<�˳��s�\��(��[_Y~+_᫆F�'L�������v�З�"O��y2���e��X�'�i��^Ǣ�4��>*ޅ^2Da0&|�mq:G�Q�=WO���(���!�.O�7.2:���u��q�a�\mD��κI�3��tf��j	-Oi�}��q��Zk"��Jn�ω�0|=��3��[�5����4[�c1�����֖+c�VqNM%�1�iP�b��;������ҟ�ae�P()��/7�hC[{A����5�׮�������I,�V�� 0���fh�"�JZ��'ћh��w��b�N��U��^R��6�͘F;�������C�X�s��C~��d�����s������k�d:�(5����[b���O�_��0*DI:Գ����E1�i����T-TI��
%�!��U��ٳ��$�p^�u��g���.�F�J�O/>;s`����+l�����}��+�B��3z���ii�q�%��}2i�x��!��B��z]�ޓ����S�9�O ���!��w���Vz)<hOɧ�c3��;3n�A��S����I6���
��f߾�~v��R_���@���U��啦�`(����ݽ�i�-���G�����d�c>�����1�F8�?sWw[��K&JsKR2�8'Ta��J�s1�j�!�Y��a	l�tF���6��Q���b#ܝ��7�R �Qv"�k~A��ñGU��(�
��9ܵ�4^k�Ƶ�G�<KF8�!4�U3@EY>.$���ҟkl�4i��J����m�vHk�Q��e�q�9�%�桡RO��M��RU��k
�yLl%��d�G�yK:�h",]������f��������05>}��SO���	 9�.e�կGo#�/���yl�H�K���A��G��� ���/�l4ljF���0w52�Q貧�٢��(�O���V�״F՟�.����a�Q�qO��%gA����p'�ŝ�Ma�b �ť�==}�Q�I���*������n����5j�t���:j�� ��%o�|�Z��S9�a�F�ՄF�K���=+���"��% x�ߢ�ϯ�++Gs�%�t{���
�klM�A��G.�CU��sɹb���',ʴ5�����|d���%c���1	�}?u�z(~x���;\�'K��|��(���E�o��|���V&�c�,D+�%��QܻE�[�uZ돯?� U����6�7Jr�mV�B�ǍMo�t<(c��7�9o����fB�%n߾��z���Xy��s���5޹;,��%Ӻ3�].�a�}�%��斺p$PX����m���yȰϖxY_ԗ(���E���3 D����p�����������	�E5���Ny�ܙ�?`��g(\EdU�6p�^O�=Pmh���8�D��A3�AB�n� ��-x��_��;�[�ft̃&��e���.��߈B�|�!po�� R���
�g������N�87�����'�<�`K�S�����iZΎ.1\�������ΐ���f�Ia��7N@ptpwf���i�^�C�!�N�3�/�yk�x���|j㌽�M�l뮳��9�x_O~��$R�Z�m��~ �	˲6_m��>MP@��>�A8x�x?�7�6��TV�saI��X��߮�ϻ�n'!N&-�!z���g�&�Pd'o@�N?�kt�:�V۱�U�8s�r϶��x��� j��8���v�:G�OL2�\iW2�	%�)�5�g�~��4��[Z�wX5�|,G�W���?�1�&�v�^�Τ��ߢ��!K���d����B�|4k	��UG^^&X{#�/��y�~:S��%w�7�l�D���B��"��&�<�?���6����h�R�\��1��^/���.�j�����bj�̳ ��pҘ9���W.N&`��ƛ������^�]���&� ����[��^}>G<�. �������V�
��u��fF���!�����U����SE2n����:�^�*��	�!r���a�R�l��E��zwB�;�j�gޚ�	��!����S&o�/�Rj6��~�����|�}������y����6�b��7^�&���|�S�I�PKnʟ��8¡^� W	
S�W��*ӧ�*Kyk)��
ձG�ʻO �PKt���+,iT��`��l������أ��N��9�ҽ��q��Z�' ��{��X�[98���!��բ7Qߌ��΀�s禳y_c��qJ� �q��y���]�LO��J�˩�ENc���s��O�M�PM�d����j����L'o�>�p����^.��U��g�}c�{1�'���y'�D����-����@Z
�'��|I��A؄�B�,��m� 6;J��d�!ۡ��zc���L�9�Q�K�@�Aa�G��$�������2^�^�B�^
���ka,�%9}W��|�{��ή'�"8���b�b_��UM�}ڷU�a��ۡÒO���ɇ�2��e`Z����TO�-K,����XGX}�*1lo":$���Tc��֫��]�"�a��S@#[-�r"��V�<{�6���[�:I��y��]���73�����݂`��M�q�z�9UvC��<�F|���+3|�A t�E��t��Y���ܦ+&��V;|Ej�|���y�\8% ;ݡH�T7� �B��WV�$mz�YF;{\�(���YvS�¬�ѿ7P(Xt�"A��]���O�8xe�bq���Q�7������X��{�m!!���:>��u�)�����m�{�'k�����޵;�b�����<�	��ss`L�{Z��lx���Z%zJ���n3kw�wb��8�]��
5�0.��5c�$�^gϳZn��'��	�"ԾK�H���9����eh��JK'.�M��Q)�	f �SJh'��?u�qF��a��|*�*96o�/� 򠎭aj:��8�9����A;�K?�p�������)�k���gKV�$ڭ&^��G�Ç�@Gy%�N�%S����Y��x��B�j6d)� ��p��+�Y�U~���|�
l�S�����E[5��K\��$��>�)�,���:(ę���	�M��f��fT'?۝��å9n�f��{PH5�Eb���qMm+��ɷ���L~S�psg^�����f����)���_�~]�5��W�?x(�y�2G�`�i3J�O�@��l}�o�Ņ��ѧp��K�N(7�M\Ƴ�J�����5���o��g![$9���;�G�3ݖ�6������z1�^��9�c�!�u?��}�h�9]�ƚ�����Z��-�.�<�Ԣ,�I)�Ϊ& U��5d��v��Sy(�4��Qn�J��j�DZF��=-�Cm�B_\����-h/z�6/ �X
�6��wT�.e���r��T�*''UYFo��"���D���z�~�xd��f�����:�tފ{�6�c}�p��8qH�y��>�q\T��T� >ՠe�sc[��
q���"����y��Z�Qq> kx:�5���\JI�ՙ~}�E}c�Cs���)�D͗4]�AU���g
��7(	���K�����J'�zt,u���e�ф��2���|��B�G�b_�P���>�U��#%?N	1M�M8�O�K_6�c�D�Z1� |�ZX��Xd�{digr{��1������Q��1�6�m���bF��<A���<�I���
�C{��̐��ó:K�]^~�=esS��&f�ۂ�L�zM�����
�	�C_5�ܓ3��t=j�����aa3gae�孵�K���<�.����3-Q~=0;NIo�o���Q�Ô�>{#����{� G�����|���o����+���l��dB>dI-B�@O��v���V�ÁI�����5�R$�� �"D�������O�Oؕ��捿�yK�*�Nq�1��o�J�JUC��9�~�� [��5=�W�M�^��2�}su��DJ.�gcB/�{��N��nQ�F�JB�%i�7gCA��5jc��u
��1��m�m��ޣG:S�Ke� �<-lTIH1��N mir)�Đ�ʇR�Dɰ�`��i��-��"�fh�D�
�!��K*�B��F�:9�#hR���JF�����,� �?#��,��>�����41Y�e� Dp�(���8��j��J�Z;K⺤��)i��e���g�����׈[�vw.ZwW=֕"�v����C�v$�/D��K�|��4VA90*M!#���C�Ғ�ԧQ��[K�w�����9tk F0�&�����A=�:F|{�Z��F���Z�}�&���o���א��j��<���� ��!���g�]�_�(lQ%Z-rS���d�mzե�#�>�����<�5��?XyAm/�m�z�TG%=�Zc&t�+H��{5C�E6��eZ)�x���Y;�k-[��7d�Q������_a�Ko�Wnm4g�9�]��!�}w�����%R��m[XCȧTjI�@QsPr������=5��c�� ���ОZ�W��|�L�R�O^p�hf��޴�zY\�(n���XOE�җ����͑b�)���S6Q�eD�+͏��b���pt���'�­�-f���.�g:���T���|�J�y�>�D���޹(G�L�.����a�"��XS���bo�z���fW�yMtթ��L"�U#��Rn�eω����l$�r 0_ E>~L~K���ž���|����@^�#�L)���
��|�>]�n�3��� ��CT7;�����I�%r��vy��as|5�ol3���m%!��P�Ҙ�`"Rҭh�bqJ�2l��,�����)����OD~J�J��
���3~��������CK��3#8�83�\D���e|ݿ2>U�MR�?gDb��O�I�?�Ǒ��V
�^��]�M��HK�<L����u��Y!զ�-���Tɨ�����|�'��<̜x�����UB������i�׍�w������ol���"��!��d�,�4��dȦCs&\ bo�f��?GϲӖ�o�9��W^����3W�s�n�"Z��4�U��]���,�8V.�VݹI�e�=��1�^п��v������~o�Fp#��Y*QZbV��;VnOש�.�c�q�x?�^~ԝ���L�ӗ<=������/E5��5:;�G��Q��#��H��OoK�x�2f��7m��B~A�[J�5(�KDL����P�A�$,�*�Oq���)$�U$��c�ԊM�Y������cD�vT��S��������{����eC�8�]��͝�)l���F�_T�K����X��h�7�l(�K���J��{�|�x_73H~-���?��쌹�Q��cW�D{�S�c�������tO�L!��!�=��c�I Z@�x�:�?��?���������p�؟Y�Gr</�s��ZQ��������BV�5�7���!W�=C$�]��i)X��ZX��Mp�r�����5�
9y������w���a���EZ��-�e�	�q�"Qz|�,x��}:%��?D=A�-ML�#�VJ3(IHc�����@/�yۑk}%���x�L�4�
��acű�o����λJT��`R|��uuU��U����ʐ���Q�
��u�r�������cp�$��|-˿+3��W��5�! �]}���1�� ���������ʯ�*��I<w���z4j���--ZB$�I��t���³���	۟�����f��P^
��|W��(�b�$j7���/q>@D�R��h�xa�?]@?��ŷ����{�o�2 �mx��~�n��\DF�WgE��Dl/���r�-Sy��{�/���>�`0��k�zK�e՞n��ڲ=� g�S��/R���Z�T�y����<� �:2��r�$�{J�δ�����x����ʞ̷7��eB�n<P��

	 y���Bj0l�= @-��eYuN^>���Δp��~�(>L�صmk[�֬}�z	K�P� 8_��jj
�8^P?�_*3�������L��>~��%Y��(PT�	#6�E�e�']������~s<ɾ.W婧��	����M&kO���b�2�$X��>�^\zN�&>f��(��\(��-��(��H�Xؤzr�I�}��G%ec҆#��C��C������\��&�f!��!>��7emL�S�T)ʥ�z,eBȧT� H�QCzod�K�����oSbfFxY�YB̬���k&'��D�y�JSOʨZ#G)�Ǉ��Tp,ݪ�1L�,(�mC��`�gWb<��?XL;���4�C��Qχ����ѭ��Ah��Ҩk���g�
�?"�:c���j/v��� !�Z�oOި^O�^��_N���q�-�ߗ�]�Y1�-v�9V�ϖ����?�W�A��#G/�N��ř_EV���\�/�62�2�2����j���id��	2N?�Q9�?�S7�s����I��R��P��y����|���k��1��e��ܔ�� �xǴ3��v�?d���͒�#�,�=~���p�	�y*U ��1�87����R�n��^�b��7��M�N���^���w�����PLxR�� P����3"�ξiʺ3�&�L//�F�
����sX������� �ڎO@���;�l$�b�_�P�����Ň��TI�)��w{!?a0v���e�C����\�X1U;|+��0Ҁ��dWh�Y��$�G�JV��6-�?]	Ƒk�V�U?^Y��3�k~���	@?	'Ζݪ��fM����)/��oH�-�V��Fx0b6,Q���U^[Y"ab�"t�l����aUR����v��d�K��F�{���^�6�?W@���DOa�Yg�j��<A��=�}OT����|�U?�C%�:%%�Y�2?ɴ���-�� �J�Z�Eg�s��n<_7�k~j�W�l�i�� g �"��O�bu�Mt�.��(�zi�ō���*�+�c��ܖbI	�q=���K�k(A���<��������̑�Ĺ��vA�]F<�덂�<���hP=��uv�͟�;;�F!��G\h�F?�ʮ�*o
U���;_+�V7N�ѽ�!�K�ao�;�S��`V#F"Z�q'Htf�C�-��I��Ƭ"�v��>�lH�`{."�gjF�P���f m�f1�{*MY�SIےJ��Sۄ������V\����S�G��u����l<( ��8���d�T�ѱF���ep���=���.x��s�oM?�O�����O���ã'��7��-k��R��YU�c*�Ƥ`�᥷1����;H��Fp1���*\
vCDeN<XTs�����k����$�-�1����jB�.��Q1F�]��$�B-/�相�:��C��g����vCiN��;�{@�/6F�6HDA@$�@��D�	6���P#���^)���`=��Ĥ�$>&���Q~��؄1�םz�J|�7����C��.�`1s9�FM��O��O���uI�̽̂{מ����ш���ׄo�������[����-t>��u�卟 iR>�}�������݂��K`T����v�5K���j���L,^�u�X&,e��A�0Z+�Y���M���>{��۱��j&�	����t�������i�i꿝z���)�Qlgߊ#w�e�򕌀P��tv����Q!C 𒡻��
�D�p�	{��r.O�^zK�a��R�Ŏ~� �$�����v���*ߦ����ԣ�����ju��3~K����%]�OVG� &;�'�@9�*�y�g�E�oe�Kg��=Y/	 k�rG_�Dq3����	-��� ��Zv��Ga��;Q�E�����N1�������h7�KL���q֧d�n\�{@��=<$?��n�I��-:):�OZ\��L������V����e�Y���ٴ����������~�Vȍ�&��e��׼QO������U֬�h��5v�2�V-�}Lx�V\�͓�5/�ȁz	�vӯ-�u�	s*��I�˨�;Y�V.-���z�3�z���c�������g���R\P ���M�Di)��\ v��n��)<�ǰl�e=��L{�؟=�	���g�%+�Z���b��Mi���J�R�}cX�΍R=Z������~X	��z�?��%�}��^��N�d��Ym�0i�-o�..��ϤJUkcX	F�|��I���[�;���"@�a?�T����|��j؞�2i�f7l���4��YL.ў�P�+7���At�xۛ�ĮB'�o��ڦ\Զ�(Wk-�c	�� w������5��\6�, [�%��XEf����G��Js���s�B��� �o���֘�����\+�u+�w>p�;�:2g����d��_a��h��s��Wn��� H}�UC��}VJa�2�;�A��g�>م �Y&��\�1H���@����"����r�7Z�wS�7�/	�xtz���d0ߩ!���j�����Գv��q���3B�����(~s����^�ujߛ�$Q�x�po���X�cB��鉸	�`��r\<��gq�����%{x_����J�J��r�8_M�.u����sru)y:n� tX�JҤ�`����8���l�Ą�t��]��r��.rL?b���P�Ț�$���ӓMn��)Cq�r�q�ے�~0��J��b:�瘖|��(�-��`* ���x��nd�2�%Wd	2ʄ������X3�b_i�z�込m�����S�B~k8F%J�I!�	n�t&X;)��A�*۩��6�ZC�{w���\�����l���Z&�&a���Xh����s��8�'�&�:u�*Uu�N�O��3e��x���Ѡ�q�&uf�/�|�N��5ͨ���x
�gF�����`8/>:{�&�ܘ�g
�����JS��K��6&�@U���r���A��֘�%�O ��G+��T�m�� ��ܯS�����ë�*Bv>���@ �Q�8��f�xK�3Xe���HvX|ퟑ����M�r�UU����N�/��}��S���?J�v�_��'�|�aEgc�}9�N�]�\��,�QY�R2�\��I���V�_����X퓩-&���B8c��u�0���4�Lw�.f�*�x'�C�Q�'3��
�3����G��~�h~f�)1xL*�,�d6���y�T����Y�ҁ��� ��g�����Y��E�UU$`�����}��S=�9g�`�f�ԁ�k�a��hg�5Y�H����������WA��ȕ��ӑ,��p���-�Ll�	�ƾ�7���>�Q%W�u  d�-�swu��Ӯ���%>e���K�fn8Y���4{��+��x~��fJ�7���;��!�A���p�F��FT@�?6#%i��X	5��T�8�D�g��^=b��O��#zWBT5����nA�]_�1�o"��e��+.���
{�})�s�x�gsUF���Dr�L��R7���_JU�ͬ�N4�:9��+e���,/�vC��^��ߋc�K�t��?�R�;��u�R�ﻵ�;��j�rU9�/E�:A`�ݝ��+{V+����m��x��I������uls�=�q��Y���"j�G �_Yt�`��F����K��֤N�(ë��"f��Z���Q��nH��D��ѡ�'���e�y5�����`����t���(~��T�ZpJ����������&�kD>&���#�z��Xrfn}�@3�!%�%ѐaגfʊ�p�h29�t�Y��ǅ|��y<|6@N`hS��R:�
�4<q��)<����<x"I�[��siDJeg���n�k�Z�_�����$��ە	����=�U-
_��1��k����S"0>P(�V�w�Ƚ����#x����"i���^�'�"��Ϛ���Ӧ��X{1>�F���O��y�x��|�
�v/C#%i�4�9?D�M�߳�A� /R��������b��ͽ���K�n	�,�fR������a���6hp�,�S��`�053*竼�^���{vҖ	| X�_�:�E;����Y���{:��a��xZĠ������1$������n���l9�֨����'��j�xA������r��&(����r���� "VQ����x��H
G̨�_��E]����;+݊�<9ю�OUUw�LW.R�zq��H��6��'`c��7�N�w3#�\w��/���'`G虁P�.��B&����=Q	��CC��*K�_��O��j2QiQ�0�{�>�}�>9꼖���	��~����#��A{�l_��r<__�u�{D�p@Y/��;���c�W�H��1�;�O� ���)�L.�!-"�sj���M���_:��dn�9����
1�A/?�3>�Ŏ	�����w�'<1|�Q�L�����'���N��)�-��yas�0̂�v�aC	�p���*�mߠ@"��_�}�nd�V�k>�O���
;���OU���>��Ukq���69׀���e+��yXN�#r����eS5oz�
1�� W{�ހj��ɖa�%e�)��Dm��8���J?s���%Ǩua���}�kFF�{xO����&�zMʕ	�e���f� O�T�
�'�W�OK�R�Z���U��C�V=ߌ��H���?LuCkDgU��F3��İ4<��-�J�踭i���D�u)�aϳ��7�P��v�wE�H��A0h�Gӷ�H���ڴ��� $x,���W�Ɂ/�͸*u�7�Eʹ�����m�XD$Ql]�,M��]JC��%�-�"9�	��V�zWmI��bd�Q͸�Y;�2>�qn��P_�_��~���/��'(��#PD�y0ǽ� l5���|��E 饹-,8{_hs^^�1�4QS�Ј�T����Lv(P�n�B�{�;��c(Y��V�6T�$v�s�c���6`9���}D�Y�PsPF�ӓN�����&*��)[n^�L������ۍ�k���%��'��ץK�ą[�(���B����m㻶w����@AFF�*R�Qu���?�㫰�Ꮪխ�GWG�� )�� ��B�YJd��7��[��b�<����G1]�*FQ��
]����ʈZu�&��u�م����)¤+�ѱq��^�L����fGz�&u
�)��EV�����?y��]E�O@��q�^UE��K���dBY��-p���!��&�p�.*KD�����&nP��~�t�u�H�C>�r
C|kzsF�Q��[���le�����G����Ð��O��P���;�n���C�Pv♦����u���ߍ��񒁽A*�22fe=�mh��΄^�C�GK��iF�mU+ ��?<��G��rl,����R��! )��ܝ'ƪ,ZJ����"D���ߢ�T� �+�s����=��������� ڞ��Mڒ�<�K�9P�i���[�cUa�Q�T�f��6�!�o�F���V&�k�T�|�Y�\�*tbe�M P�.� i:�yH�V���o-ӫ�5���W�-s�u���w_�'��8�u�bi^b]��T��c�W��@�a�ؒc�Һ	6�M��\E�A=�*���M�^Y�%n��|{�ڋ�GB�t^��:ؚ=�n���LXi.�Q�3����E�o�B��s����ʂ�n��5cl����t���e��N�����[O����E�ƺ���ɠ���p[n͚�h���;�z{�C=�fA|��w|�r�`��u��c���x5������:?}cŭ�yysʿ�[�Ǿ#z��l8�Ђ��[|H>�hE�fTG��\wcUrO���.�O�Jr0��k�G�!�At�0Y*@�*w@j^�p���9Lt5��x��'�Rg��k��/����y�j��%EB~"�r@��0�q��M��~�y�Y`y�[Һ)k��mTOlo9sF��`���������4t�Є,KQ�O��(뤔@��b)u�Vۥ�3s�[#\ϣx�����/��,��q�u[S�2����VI�O�%º5mt�W$\��_�]La�V8���ha�JJ}G�M��*��@�2kx�y���G��F���_,��@q�Sd1>t{���	9n��Ι.75i9Y�W^j\w�/Dl�Ea��R"�������Ì�}n�&��M���N9j��"~9�c@�F,��p��3��^�^��K%��B���;"��HBkN��̏��3���}�����0t���lY���iU|VPZ����[� 3*���fQ���
I��c�t.��7������s��<�'�<yR���GPb�?�]���D���nkbϗo�pTmB��1��J��;�J>L?���\�T�����)�J����t���U��@I�l&`�.#/��1�7��+Y+���ƦV���f�9�8��9�G�Α|� �d�o|��P�RVj�����;C�tW��9S*�Y�'���j�S�'��Ԥ��9i�Vs�Єmp4�K�����h�}{NTooZ��O�P~~,��?kEFb��k-O�}�����{����U��.Y.�	��.]�E�Ѭ�5V��O�T�����1aci�%p���A}�-��l��A[�Xh
�T���ߒ���F^̲O@[&K;I:�Ti=f�S��R
U��hy
l��)�}����.��fV_�^����Y���t�	�	.����H�@����A�;��4�.Ao��iv�k����Q�V�9�uW͒ǝ���ݠeז?dl��3�P��r "�q&�++T
�j?li�����<�U�b�G��X��QB
q�>sbI��o�O��O�'��� o�v\x���âR����К����I�|3�6�|NL�F����`)*�� S%[J��h��G�U�K�� O@�K�b��J���a"ǃ�}�=�
x�ƿE�� �b�����Z� �T��Ҵ�b��k��U�8�{��	e�2�"�5�'��"����4!����?�����*�,�fI'�R1ꕦ𖗇�,��Ԛm��1T;Tf��o��X��{Ꙙ*�\��Ctֺi�P�;�=����M�	���Еo��/Zb��7@픶��@�3[_�uY�&M9M�%<S����h��Z5Z���&e���A�t��y�=���2������E;Y�؟�c��R4�ǍU�(��;�\x�I�ut�X�%��_�t���+��>�Y�c�oW��Y�d��W�V�{���(�Ե13�h\lYz=V�w��&���}�ZC���ӽ�ݶk�������o| ֆD/�_�����y8��?=�=�"$V����)�t���2kĊc�kS�\64�V�ly��.N7��kN�O�/F�f+g�����?��w�f�����2��u�hs�/�Ч.+qEm��^+��n�8ݽ�x�,�ŕ���kK���c��1m���K2�h6���סl�����	��b�88c������I�X&C�Y�ˏҔy'�����{�v���.��#?ߏ��dN�����M���v{�p� O��P�{�9쓱GI�}��|��>�L���Y��m�JI�
r
�O^ͤѤ�t|y�%ΪĊ���\�?Ĵ_G��"�0q�;I�9�ۯJ�jx<6P�+�*�U�^"�x���/���]ͩFK&�愇fʩ�A� ����f���#G�v�{$��䓑��K�%a~p�%����#cU\�nHm�N��B�ϕ�}ڊ�Wo��n3�BX6Zc��qk84�E�p����Z�*�!g���G<�wy!zӰ7 ֫>S=YS��р�n��ju�������mV�
[z�x�R����;TJ����!�ؼ� �gX��b!:R��\��ھ����wId�x����B��z.+(����Ѵg�7�̜��.�ڔ�k��k�N�UN�D�>	���x�8���pBE^��^�N���34Z6>/t%��X�V��[g���MO���c�`|�++����|��@��ױ�m��\3���D��z����-�B�d)��Qw�Ht<<ӧ.��7a���i-��~t��HNQs��Q�˴����}*��Xlc�	�9f���Rj؃c�J�o �gt㊘'�4Q�����Kg6S-�ݙ��p�C0KP�o��{�4�2Kd	���й�%�H&(���i�V��Vg�X���f�G�J����`?{3�$H���<x޶��~�| ��<�3�a͠1B���	��������,%ŋ���`CԮ�z�"��a.)D��'
?Gpe�W�xHV)�&��$����~m�r �8�.�*�+�)+.�O�����e�d&�K���n�!Nݕ"һ"d�a/����r��_(x~a�Ǚ`ĖlfT�S�MH/'*&�#���]�mf� &�QI�tE�FjkL�]W��V����P�R�7����{�oJ>�W���ԥ�Y�	�r�!��ze�I
bJ�߱Ę��ieYɄ�����(�>G��h]�	ɍ�KɭW�S�)����q<��m���K#�t!ߐ��y�8�4��_S�p��j��52�J7�z��4n�p�S�l]<`J�Kڍ�K/�A�<����!��İRG��8T�hs�0�6�s���s�9;��t����3vE��hEZ��F� ��F�p�Fm���.[-\���������R�P�&�H�������^�5��_ͳ�F�P,��	w?/~u�g�֪Mw��>{9a�ctz3^���٫7�w���~���Z#4��f����r)1�	{���X�~<�Z�_���Ũ?D<k��Df��h�ݮ�l��j���n�'�io|�4�.�#��B�y��&�k���H� ������I��'?��Z�X��6���[�p�u���W�*��_%�T6@����Jv��-`�������u�7p���ne��6a��R��o���:ժ�eWk*�V�N�񩤳�VE<mkP��7�jhm�X8�-W��V�y	���-���
��4Q�Q� _o&��y�X�/ҙ�(�-�Ig���@��_=5�W?��@k�8ieM���z�b���ā�6�Oj4o }�[MlTT'9��7 ���E�ڴ聗)O�?���@V���?��sW��~����;�;0+�.��KG�*�m�N��v��=����_�O��Ϫ�#�g����kD��YA@���W_F�1�W��M�-)�>��7����O+���E����ԶS��ob�&ګ�������& ]����h*�s5���Yo��O2��묌��)��A�Oٓ��'�B�-!��A]�I�a�E����w�r+u���G'CCyDi��>�+)R�
�+��*N�2���5i��䂝Nv�ObIq�b��\�r��M�;�Z��p$��Z�C .��5����{U����;�����і�5�v�7��.5�x�b��g��7��J�J{)�3���{q?Pě�DX"F^�h��O����Uӗȅ�����;�R�B2�|:v����+I�����W��Eʸ�M��X��k��ng�ˎ�=!���v�c��l�������)tܞ�j���t����ώ&J��c�H����w���`���ٲ�q�Tv�A  N�����n�;sGl����W@3S?�[�On�>-+���}u�&�u�v��u�$n�zBi�{�T9�n_I�w��m�lv
�rdLeʿ�?)��9�E�m/f�C�a��>���T�[*z��A�ُ� N�w_����I������܀��9�_���XT�y��d�%r�3���&Mϯ��/�� �3��T��Gڏڧ )Q��:
�W=��s$A�?��wDe��&l����GU�+��� �J���O�}o�D������J�9s*oC~B�ͼ�c�����,��o|�u�q�4��MW�#�)P3k�>8��<-) �%��������?�%�D��8�V2^n�B~2J��Qn,����M��:�p~���ݑm�bf�EL����E�_�BsO��-<t?Y�wm��^^��wX�x?+XaҌ;j>����yL�5śS���I�\|�m�GS��@�l�.8h�v3k��~�g�u��g�9�j��fV<�v���L����)VB�Ж�V�Ǘ.%b'|=�h�� ��F���L���j�Or�p���*^ʣ^���Q��0\`��Eb_[�dC��|o�)L;�/(��p��(�n��������Uo�z�f�P��|u�c���m��l�V_�s�(�CK�'���r���~/W��'ԡa�%AU��`$'�j}4�e(�a@%��4�i���?����g�`)��2�ү?E�?G� $!���]�*��qyy=���Z�o�z�������N��S������4B�\�V�s���fI�ĵ)�ÕBA:C�3�t8Ox����&��LK�ag�G���k�ߜ��mU�J��;W�(��l���-�4���&紶��e˸t����WAG>�c-��rU���!G�~i"1�p���:%�Rd6TE�wm�ݪ]T°����4�������Ò{�Q}�Ռ_f�b����J<�8O�{���G]�m��!P�JnK��A
W�O赗��1#Ǝ�x+�T����z[�=
3�N��w�`э��L���+��,)}���w�YP�8)��S����5�������6�E�NV�]���r8*�hR�XɃd�� ^�8I���J��耵�͢zY\��ҼS�
\_: ���Pk�P�Ϯ���g�-,�@�3��7�w���`��8��}1~��)���QqNTk?_<��ǜ�Z�!b�5�־x٢-IHoS�p���O���t��M[�zf0�[���g�-�ե]�aM)�U\d�&����_��F���~�1!+Kd�-�#PYy���1�T.��c�{���I���'����<^�	W�5h�+�ǅ�9^���]��K'�D�����HTaOZ����L��+����8�toh_�md],��AʮY������ZZ�
�x�/�E���a��
�:����v'mǛP��+{��W����;����Oed&V:�{b}d*��&x4��̶?!.��o�H�7��uߩ�T�<<�r�'��=�@C�?j�w��b& ��~ŧ�p�!Я`X+NǞs{��$!�疞�v�g)\s~Y���1Hv��Ta�e����>��_6g��1�z�?�~JG�)q&K���E����C�v�� )Np�|�3L���=�T�<���e���Y2�J�e���u_Ź1T�7b')r��s�D֨��߸F��M}8d�j?>\sn>�Ԝ}Y��d��)l����$����e�oO�U�ڭ���U{K���HTG�j�� L�XW��.�'( ��vA �9N�����FK9��2:F��[F;�[5IJ�d�1eUH�WD\O�r�Z3��_�$�f�)6����8�Z�M]GĔ{�9w��Yx�rW��\�D���B*�����"�h�������?yZ�-��b(�R��旘�>b����p��|�#��(.$��*O,V�8���a���ƈ�G�sRI'U��BU��
�$}�m"ps�?��y�7��@�e�N��·��Hw������f?ᓁgě���d24�/��ѻ�W7�ξ�V�?���g
K��\�qE	Q�sVm�o)/���r��p�O|�����J��Z^8LMF��#jE�.�[@��u�_(Y�^��a쬋f�p������<WR�dTg��|�5���#��O���&�Ş���z� |��o��q��#������p����	^����T$ଛ�F��K;�N��0`��q튳qb���Q�2,��h8f��R^���_d\hVjk<�'K�Ԭ�� ,���/��b��3��5	�<�l�^� ��t��a�Z�Zi���W~n���{�P{�3".s�s�7���6��B]utm�Z����w�EV鋥j�Fc�{_�n~��ZS֡�N~��Hc�f';�f�g��뜏�9�=�*�oB�yI�\A��a�B}����ݶ��׿~uGQ`	mx۵������?i���w��e���9���ak�#�;��V3���է��G>1�3�15CZ	 $R:L�X�7�}������aLVA����j�ƥ�9c+�Ҡ�i��t�[��RK�s��֋٦�A1���-1�[�8G9��G9\fg�[H��秙ɒ�%m�S��+kZ�M��B�QET�a�
�Cʰ�Y�?��!��].,�����f�q鼇���?�-��B��a|8w�dp���ݮqv��ka�8d�(�d�"5uF���#m��JB�����ݗ�]\c��-���$5!f�T%�^�o*֮La����/Tu�UW����9����r�S���J��bi+��f�O�#�B�@�fvb��X�[4���Ѵ�� J&�2ai�����N��%פ�����%ǻ�bԚ����_\N�Fz�r��S#�^*��θ	���L�����,�<q;��-4X�����ac��̥�L�UO��ߜ8a����$\�^=���H�[i��}R2��-VȚ�P���)��j���AB�����k�m�F.Im�����׎����5]�&�ܕ-�����5<�7Yv�t�]�+�T ��W�$�{�ht�k���oI��l%����l�����>wb���(�+����;�!�$c%W���Z�w���߇�.���n���Ɔk�QN�SI��r��9eGR��� u��B�ij�X��]�� YC
�/7�8B�^�i���A&����U4�����;��d����`�����Y[��g���~W�5-+$u���166�w��+�.�	�L O�'��ӕ~���P305X��%�T݆�$C�Y�wï��f��O>O�g��t�>�R4��3Û�v�g���b����Tk��|۸�,����������fl���,��>�D�b ) Vk�F1/��+�6Mg\��툠���5�
f�E�ָF�.[�4��7���=ȿ�+a�?�6�9�.g��1�;�>w��K���+:��W:0"Q��6o�<�pǻK����������B��"��@�^��I�1ȑR��A�W�8
�
>vG���	T?�� ���7 Gv�ӧm��{�K�.7���?��≢�E_�˧�.6+���@g�$�JRB�E�ɲ�0	�N֏U��<}� >ֶS�Y!~�#Y:\#"@�جsYwB�8�P�*Nꛆ��Fz{:P�o��T������(	KiF9D��2� �� ���|�"�ԇ G�1m��A����� ���c$n��6�**NO��۳o��J΃�<RgU�v*��Ƒ9 �wf�n��g�V�J��[�I��C���o����7ʸP3��!�Ђw;~E�2��7�wd:�c� ��)Z�w]��R%�qI��'��*�6�NB��קKq��D�q�+fV�q�����p�ջ1���o	�R�?�3���֏O��JU�� ���rr������y$��T.P��B#�a��[��d�In4b>[_�1��o!�W�3��2*ͧ� �hqIh��-.�k[����v Bvb��=�h}(E*W8w<���iHY-Z_�U��Z�Iɓ��J�L'{����<uvIW��
��V��<V6��#�0�� �HHeuzzBD�1=�ots�_Y��ޫyfI©И����$[׆L�OR̳4R��*�C�]�oJ��*��E�d���x�����:��	���҅ܭ��q՝ᵖ�?�t
���{6�n?`u�9)�a_VL锺�	V_�0��3�[�&�WO,��h?�<+=0��d��g�u�6%�A\��3�ݛu4�cX_U�4b�5�wT�T4����λ�Si�%Abv{�͕ޚ?f|asm}���-f��)�f$�����T��-���w��.�^{�l�>/4�����exp�^���!��o�U��?u<-՛��}��<�K�%����><�*Wjju�v-,�
�e�T�[����U��U�-kw����*<&�s���Q6R��ӎ�����VbDz�;���ś6��8�K�x�	&�&e-�[�`�7gs	��q�7MNd5C��e���b�!���K6y�� ;���7����9�,�"q�ߋ�xv;�Vܴ��6G�/Szp�)Ձ2�1�~��T�5C��:r��<��$*@���b�����9�!�;]ES�u����9�����'��n4N�9��r�_6\;&�X��V�኷A��\�>� GW;�/���"ƨReY��z�*�v?Ϩ(�9�+�H�� �w@לּ�#��a�\�[l�^�+�� ������L�KVȷ�T��L�&�:�Ԑ��c;Apa�5�w3_�R���'TɃ�X �\�n8\qGE=Xfj@0׼q5�ۉ�ܖ�]�1��>)N}�����\i�`(wi��$��,K���ؗY����kt�UU)�&So�U|m	`5l�w�Ζ����f�}�d; �ҿ���'��BՊMڲ����������D�����������������l�ɫ�73&��ڼ�/������7��p��t���ړ0O������q��?���ds�;n'�,��R}�`F;��!�v$~T����!�T�ҔlTi��I*��ǧɿR�1cm���J��6�;W.��;F�x���N~A>�B�9
E����P yOI.���n�F�����Yj��%k+�g���z���]��� D���R�|���V�u��	���yt&�݄�ʾ�'�7�l���)���"-c�U~� $#�*� ���\��������
٬0s�)_zG����P�m��f�c!*�ϸ�d)�����ɫ��������3�&�7 ����e#T+�(j��~ˍ��@/��<�G�	zq��8�xTϋ�����R�{�g}3�U�.��Ig6��Y��>fp�q�@������<���~���(�>���� ���b���s}Z/��OC¸�f��o��Ǫ���Hϛ��	��܄�ゴ�S-W��M��n``�
��s�0!1 $7� ���Ү�?�@�R7^���U�������)��^΄0�?-��NϾf�O־��a��˒3�S��s1��KU�h#9�2�c�+��_q���qUʪJ���{��tq
��=q���f�V}��^xp����}��ƶo�m�j��(�i��8Trb	#�
���1&��'l���J���|�K��;�U�;��+�����W(�b�W��Qa�.�n�P+���MZ<�d���H�d�r+�h�uN���B�u���qx.�@�ѹ��dk����B�#>��car� �g�`�����*^�����V�A��/�û7��iɸ�a)b��l�r.�
֌g���M=�p�-� ��8��^b��aR���a����u|+%/�5-u��Q��ϊ�%K���\�G�PR�`@W�^��ђ��|E�?����iYԱum� ��E{4Xp����?pTy��!^�N�`�oP��"+���J˾�&S��:z�������D���R>h^�p&V�����ȧ5��>c8ߋ��>c��еn{u�& �KyS3r��NGC�ޞ����o1-7�ކ؇�K��Q��`�������iC�>������e���#�nǵ�.��d�k�(��0;�6�������B��Z�Gd�҄��|����;lR�ȑQ]�D���$���]z>��K��g�'�kp'�(o%O��V��F,*����D���m�{l+sv�)����o�1����p��(\`v]%��D�_��v4UaUv3�̆�������\��dN'�b�b�͵�Dt�8��[e���G�-{���Զ��o��%�|��h���K��:dI�εo�-��z�����ы��2��1?"�:F��R]3�A.٣�{���O���K�6~m��x%�ʨ=c��1��y�:��l�}�f�ώzUH��y�U��96�}b~�0�5W]�_�,�y{� 3�U�ɷ]ӳ�z���(��o�ّ��TT;����\��:Y���4�հk\�|��g_��)���\uJ$d�R��Z��Z�ژ-mЫ�R�^�G�Be�i�4���(�,��H������i>��jj�6]��bH_�Vc4ɽ�	Vw��EN|+뭮�#H�N�
k������.{Mk�};�1E�_��ْ���i�ui{W-�eo����9�^�7>�هE\��K'�ӟ��L:�,����uO�1��,s�ҝ��;��/r�_�Y��ͼ[���y`⾫)v[��� 'u�DuUa�\r`�Uh�|��U؇�9��2!�ʒK��C�|SKZ�0������V�:*�ndL�
�
ʗ�(}V٨Jy�Ձ�D�_�S���g��g��`��[�y��� �������NYY׬�26L����VGj��k:��
q�%��UE�/,Ū|��(Jk}���8��ʱE ��t�XS�aN���]z~�
��Z�����4"�G6ΰF�w6S��Y'�ZЅ9�����%����&b	�ǔM�R@�ĕ�&�mQf5�xR-�ߕ��í��.�c������
�F��xE��rR�C��B�f]��U\�?}8Oc5l@:�kB�g�*>�-^�������D�<�l��C+��;}b�w��Óf����JG�j��9����X̎�7@EȀp�|��ZJ�����P����׹xew��s;z�^<V�R���T4[�l�(!B�"e��0Ck�EZ$]�y�I!��#�>�W������w~ݔ�~��A �oo���?@�o�� �lĞσ�}����*��fE!Bc�;��L��>�=�=0���d׀��YR������xC%%uTϵ�Y�n���[@�bP&o��C��O��@��?+t̙N�{��G�S�/]��:�4�M���~��ǫ/I0��7@��U]�5�-vo����Ơ�3~���^ca�1�;V�/%!��4� "���e?��|=a�G���˷u�5mS����{��29��-y���#��I�=�@mx�]�	uv�Δ��wR�
�F���~������|�����'�KU�G�4w$σ��T�����ۡ]v��}�����x�T�D44(�V�t�\C_���Ftj�yMv.p��ax�����6ɚe��jl䕪��[/WW"�q�R�����.���X�x��JۍH�$�V@����d�W)�f�ؿ��Y,I�ex��N�5u�������"� ���}2z�,&��J�^T�]�Į�uvD@�B`\�� 1��L�Վ��r������o����� Gׇ�	9�2�s�+?��-�?�������El-K����u45�1y=80)�P�JJw�����`��A�_���T��A&0s��'3VT�r��3��(ֺ�i]}�TJF;`��i2��?O+�ӥy��VI�Q�6�(����Cc2�������߿`��TZ�x�1֩,Hof��/��nj۳��Y��u20'!PV�9֔�Z���a�!����ض�	���v\�\�4\�?�:7(���#�QO	<a��ɝBa��]9Xf܄�j�����>�HZCp�N����b[`���)��*;̯M�_`5wo=�l�]�<̆�WT1�mpu�b��Å��N�ɑ #����%Z!M�Y�M��~,��MQ���7��1�Eȑ	��Q@{֤D�����脺���"2/�|�C��G{2҆1D��C6u�RyJΉ���썶I,$V�ڎ��-)�����9��OR����J$g�F�ǰ�u��졈�?5�?�4q�Dw&"��wV�]�5�ˏ	��Qp���ё�+5;�I��|�>\�jݗ�A��zjA-G�߅g�+;(+lO�3��`�����E0Ͳ�Y°I�/}�6���d���?�t�7[��\���;���JX��Ɂ7C��M���*0�j�>i����g~�P�xT��>	">���O>�G<��9�i��D8l�_�0���g����11İ��YT��Fg���C隭"G#��B�O�)�&	��=���}���S�ų��խڶ���w�A`Z�%��h|�Y$��R@�t��\q�wbs�����V��@�X���U�Ҭ�o�F��p�FoorF����D7��5�,�.��
�
1J�4���8��SH�=�]v���f�.��+�:�r�}7iУ*�b���������ӱ0s�L@�P�&�MQ\��]S���=]%v���w��o�L�v������80�kw��ٯ�n��h�8=-�.�k0{2A�Z�?�ǩA�h Aǧ�Xf(e�u���Ha��'�]��$�h�v(�,�zDpb|x�vڤn���y�<�hUK7;Nj�N[2�j�0ŖpFbp��'�z`�(J�A����: �C)�t�S��PQz=�)�MbKO�gQ�05I�XZ�	|_���Ku���.L�x*7�?uD�\	%P��$�h{�X���_��(��/y�O#���&��ڗb!OIm ���+��ɐ�����ρ��o��'�'0,=���3��Z9$j��jbeHV��B�8R|&W��\�)Ol=C�����H�k�����^����j���9@����P��D��-��z���ɴ8�k?��IW}�؜�34��`E�_�S�0�t��ae�)G.���8}�{��7ܹ�+��rWD�;��Λ��i�ȍ��rq�����m���~m͆�*��N����u��A��$U��|�m����R	(d���!p[a���B����2���"����I�������7y}c��!N&q�Y3a^c�h�|mD�?D5����\*��B!�4y���9��� �Uoj����t����`�A��Ў1���PVT�{UV�EN�/K���U�����~���>4���T�4a$_��M`B$Ee(-[�l�j��'t���uewW*C��6�ra�P�p�$:6���T%$F
i��/?�IU2�އ'�����_iC=R'c���"8ۨ�[�4���C@a`l��xs�u���¥+!ʑ��3��e%�+���<o�d��zFِ'z�ͅ��$`�9̱4a��� �F*6E�t�U����v��t�z52*����q��YLzh�ـ�b�P��yQ��ɟ�e`nܙQ ��r�M�������FK����2~�kq��O��ܯ�����6r�"����tOb"���¾K�RՏ|��z�>}o�4.��z��Kc�ٴ��G���v/�5u����ݶ����aŕc ��uqq!�\U� ���6Ao���;MuV�{����ܢߨY��4�:���[�����5���h�ǣ]O��z�l��4�o�֘�t듳�&�e�����1����эޱ-���Y�l�LI�9"�d'�_e����YYɠ�3U\�}�:�_��߂-ޯ/�KDZo�Ō,-���z+��d���z�۶�"�TB9C�'Hز��̊RU9f����V˽W�2G�ܭF5y�g��� aa��*��5��\,eJr��� 6��*~���%!�����W��}H��^g����7��顸W>�B��̓1�M�|^�e�%��E%a;/��$���׺��v�`×J�K5��N��VlTL�3�
��ݟ�>���O��R#����|vWCA�()Rq	UrJ�K��Z#�k��?J��z���1�؞WeD�ǽ�A	�1I聺��R�z����m�WV��8T�@5^���b��g�]]b�����|���Mi�O:
�4}{pG^�U�����m'�O��E!��䞸.ul��Cd���9���`6�Ų�QO����Ц��U6�U�B��x��w�^���hx�a<�1Y#pWQK�A-���-�􄿵=]Z^��� F
�\��bv<�{��ۭ��ٻ��:5c6�����>��;�D!je4A	�����#�
d�P	k�y���4{��gj��dO�%#�ea������Y �����q�D�A3m����Ϣ1M���X	z�x��)W4E�>�*ڑB�Q�&����%�����f\9�������
!�ߛ�C4,����:��e����z,��"F�_1��������Wٯ���"_�[#=���O��Y�
<1Ir�FEi^��W���(����a��g�4sYg�w����o��2����P-��_��k���h*�\��%/R���{�/�	�қ��}�]���l�,
�����ۣ�7@2i���UF�,�?�o���j�T�+����h����Y�5�V�̼dL?=w�ם����;���l7wO;�t���u�`pWO��e����T��];�#=U58�`���
S�����dR�w�x#�u(���P�g�jf�Z��`��q�W�����Uu~|�/?,~5ϔ���=��
�/�啑����NT:y �����Kp�ףkg��}����i�-X���Ovp�]��b/���@��T�;�����' �"�c�Ŝ���)���,zZ���VVV^��Kk	m\�ԏHJ���5��N(�Wo ��ʏ(��i�}]�Y����w�^Kw\��?��ͯHnJ<u���xY�����{C�>U�G(����)^'*s$,cd��$�P3�<C��*DJ)��,X�����K��H$ֹ��<,���])��b�x�ҪU�A��'�{�:�X1z�!��:}�����ȳ���OC:�A,^x.��p:��[��'����tϩ��[j�Kݡm� 73y�d�����((��jL���N�6�~ίp��/,.��K���aU2_9���V��"/�B��񴲹Wө,�[+K�85��U���ܳ�f]�X�Y�����,]_!&�$�pe̟�Z�E��0<7y��o,�֒r��/V�%�7��_R��?��/�6a,	�\��,qƟ�$��y��D���<:�Hܥ�Ң|�;4$!�ۢg!NM[��"��Ǻ0�v�0��l�"|�K����®���t7��֐�����A~򔢉�yH:�C����}�A�'N�(̴�zC�Sy���u����k�\&�!~淮�\�%�j?�4�^P99�)�*�(������]}��J�T��O\o�Re���⒰ ����yB�� �Pv��8��� �V�C+����Ȯ��_,���]_�GP��y ��Z���sx�+K̜��%�c3�(u�>FQ=��l��C�E<q�"Z/f��V�=:T*?(%1h��pHq���

R*�(B�d��8fg/+X�!�����*�p�pU�� +�o ,��g<b��jM��[��aR}��i��뙐����m Cf�Er���/������I�}9)�$�4��e�u6��?���}Al]�qᗣ�+	̂{�tC�����H��b5Z�����p�'n�Lmт	��P�o��$�p9��SӾ�?�}������(��%����\���h���ɛ�O�ۄ�	�^=�����i�8�g��/�Bg�|M�)C��^���4+�{���*
��Z����^�A�����¥A�K �/��ŉ��&�lO�B�ds��ǝ����^��)�rv�TF{� N܎y�t�ʿ�U���.a}�搁�S���M��Y{X�n���C��ŌҿB�0�����LX�=�\&��+}��,C&������_���I�TȀ����ў*�ܔ�D��ĥlА ��,�ZP�T�AT�Rkѕ�>�~A��|9[�*/�����χjwW�Q��e�>�
�+�M���И��4E���+��f�#��gqVr�{H ���*�+{/
Ł��X��&0��s�bEJ:S�(i�_/�@+.�SL'�ڏ�e|�܂	At#�o����1��}mx����x<�6DK]M�Dr�J(y;�$亼/p��է�r���Jw�	�^M��BMTU�LzM������	����>b�o�9�p�y��Rx�@�{]g���cY<\-:ZVl��3���������{w�Ĕ�N�����`�C�
��O�%nLb�������Վ��w��L%����LGU%y�+�J�,t��@�89T(w֎�J�OP[[���3dT-t!����9ھ��e(��j��������טy��J�fĈϜ��"�Jz�.�2�mN�c�'�7�,`(gr��g���|�Xu�SL�V�����k�Uf�gd*���L1̂>t��m� �i'0S�gHG�S�_~��e�	�ܠ�#{���Dn���<�����(����`�i/=c����Z� �Cn6뻛ϋ��B��7�Sk���M�̄�iMg�~��^�USsNEeaQ��H��6�ZVi@�r�i$���pH��8���#��Z!�	�=� �����[;ɧ�83�
��ǊO�{9h�ZsN��[_���G�l%��x�ā}J��\͋�fPV��p%�`K�;�ƅS���a~5����+�+�~Nt�k�� ��P2���M��΅�H��nA�-��KP?S%�c�d�F2�rg�-�Cs4�8���ITꐎ���ҫ�%7�8��X�A����M�1�JL�'��l6+!ս|�����e��.��,(�Q�Ub�`&B��M����eɡ�F�r��m�}w����Ҿ���)t�Vlr�,Q�1�;򺦚M�����D*�����IB����!'u ;g���-@¢G2[<���Q���=�l��@�Pu�}O��-XR)a���t�,�F��S���ܒ�>�8
rM>���j��;/L��/�F�\�'�J֬��~��Rkí�	�3������bST�|I��+P�cZ�G�Ĺx�zUH�g볽���a+���^cXm��ǝ��f�4`�Cӭ��9Xh�vL�ǀ�Q��܄2���-��>�I��4uX��v��W�X�_����ߟ��.���ү���g�@ո��x?a�xi���k]J��w/��'��̌H��~������1o��^��j�]�^�w����ݲ���*۴�*��Q%�����o��e��v�f�� QЯY�o�e W�qL��Ow��$�O�,7�suA �P1��4���%dђ���Qi:#�S1./ [f�Kyw��J�өg��}��G��w3\�9ծ�6�\���sg�Ӵ���C��$��� �����.C ��%���n������9y����e���U�]�U������0H�����=vT��ʕyOk{�	��m��������Fѹ�G�yH�8}N�=u�xO�C�a��Y@[�̕��,`:��QlM�e��n��S��݃\@���6���s*N��v���m����&�%A�/Pe�_v?�ch�j۫��h�	;�*�ȿ�Xm,����(�����9��(J�j��%O�E,ݜ�w�������ʣ-��#����Jq��?�ᄩ��]�a5��?!�]�&������R���
�c��Cs��ަ���~���ƅ������cqrL��U�hs
و�4�,�5��\��a���M��f{!�)T1����?�%��Դ����l��~�<���윘�κ���̡�䛔���;`�;Z� �4ԟ+ e7�і	$2�c�g��ٸD,������u�����K������HwJEB��;������ܻ�|w��`�0%R�	*j�>�����O�E�C�O�����6�'���e������1��|�#�n�CU���U���Go6?O
��C�T�����nԴ�[l`-%6!����yvXX��fr$�G���Ɖ�a�Q�/�x:��L�O�5?�$�J�aC�n�e�'�z��^��iv;�c�־��QI��+m��sf�W>�'}k�Ij�ߛ�7���k�.E�p�y�j_V�Bj�\�W���UWg����l�Y��W&?�a	�=��K?sM����A��-A|��a�F�.ʜ_��1���=��C����R{��?�+.�0�Һ�ɉq�:R)�[��5SF|s�8^�v���y3��͒�l����v<��S��Z��r�E	��8E�$u���U2֎4�!��\�m3K��Y����#x�S�W�����1!����БW�0-�e#Bϫ�⦄���tQ^P���߃��[�&G9U��I-hW���ڨ��+�R����'|�Ӱ5���5��`drJ���~��w ��V&f�!����ֶ�9��R�,ĉ�����N����sv�Rs��Q'}C����X��嬖�5tM����&��	�K�RG{$����gu+�+L)�i��ss�G�{~�����oEmv;A�@�K{������OFe��yRA�x�� �M) \ ܠ�7�t�O7�pu5Jk�2��'�sG���&��&M�2��`Ә��!K��|�r���[���"��ˡ04�p�X� ���q+;�}��[^�2�T�	�_M?�c����g!ѧO؀GPv�� 
*?U:&P��ꖶ
�/�R*Z�I���/�,n��j�a��6�;ʤ���t6l��"5}�[���틩0v1������HN~��9�V�^�o���˪�m˕��rk��+��5�mq�(i�)�n^U�;��'6���$6����z�b=���?��!�sJ~�#�7��3I*3��lM���?�p����1���+U�k�;��m�����	(��V?.�Bp$$�<5���+�qS�ǢCWLj#��龫X`U	+��=^˭���l�+�v�#�]0�4���XHbj��u��>�l����2`�k�n�]�[p��2�I�l�k8�=�}wN3dok##j�	����_ܒ����0+�
 �%̹�x�V��:��R�*�d���R�M��{��4b�Z��j\U�X���P�S�F����7��|fiQY�
l�����td��3##�c!��Ä��<�2V�X�?�4~���Zq?>��'��M���'
�m�xϢo�:
%�̿�n�=�����d6�ͨڢ)ޜ��nGxJ��zV����=��\s�a�����9Z�/׳���X���}����u�����43U<Qp���8���O���}/�A���5Y��nGnkxL�A7
�?�Cs�e)�|�A�����#Eo C�����	~Y	<���G�ӯ�YA�T�+���Y�c+zG�r��.� [p�d����?O�=<4�!Q��c/�f��m����z�5m&���C��mJ�~�fK��niu�\JY�h�B�dpU�6���	g�cτA��t��0�7��#8Ş)-��H��u��q����;��D��Q��et�Ԩ�(&*1#+|�9//��2Ѯ_�v�|[�4���^�~Y���V(ʄ��j�7�d�U�����9�h�7�6fy6���z�P*��b���ޡ6�v�aU��(d(6��Sncz�h������&��-1��w]q]ao �|nմ"�ٙ4fE�Ze���I�W}y|��,k?��g78O4׾Z]�6N|������ � Z��{3�@�$eI�iY�L;3Ƹ����wB�xR��AT������;�^Z������W�H�;���[5k~;I����޶�_���|��HZŝ2�Y�[_���Fx�w���}��e���<E��Z�s�Nve޸�yBX7d&@���}�-���"�Vi�Gia��.�W7_@|�{�� ��Ϧ����2������fI���<�d䜬h��Vj��0��N}��$�����2��1�Kv��c��
S���z�*y�y<�V�_��>�IDrc�aA��,��x4!L�
2s ��g�������FN/���#9/�|���&{�����!�v���Q|��59�_���������jo�;�6~0��;֓ۛ%�V��Q�p����ٙ���Je��Rf3pV�!1A 1�������{ xwy�����ٺ���??d^�+�)+_[F��H����%�Xx���O�ĝH`4RL��4�y��S��q��� �_��m���̷��a�(��8���X�H�CZ�r(��P|.}�4�R����8r`��$�dLA�p�T���n��T�*�֚������͝ɫn���*����Hijr�6���,��PU6zd��Ө&�~��.��;����U�@#ִI͌}zmci*Җ�n��?Z�w	<��kI��q�:"o�vss���䦋W�'乸��ԡ��EE%Eq9%aSݞ;�Y�;�u�q8�]��@!#��}�S}��{ҧ��-7RD��5�b�*ӧ�o�r��|ڡ�(�&�)���Gq�;��*Ż{�qċ�E�b������j9��C-d���/�~�@_fSTTfm���{��C5Mk�YOsI���Y��&���t��׮`���a�5F�*݃�4�_���8T�_�m0X��3�dЖ�G����R�! n�/�z��6%�"Żo�ڥ�jb${�;�ӟ�Y��f�K��l=��ڔ�"��	h�C&^ViZd�("��nhƤ�����p�g>�e^ڸ��m�Z�>��7�{&Q���g7�8�����~�'�����$�Ź���<�'R�>���g6RH]D_��� v��>u@-;5��������H�O{�� g� ���?{t�s��7����������� kT��,��>tl��hatj��b���?z��o��E5�S������b:4�c���j���QXwY"���~/�֞:x~��XA�~�(��L��*��x���+��R݊d�����&'�$�B��M���-�j����Y '�S��c,dt������l��]��T�Ĥ���[6^B���92���^�`����4�_�5���E_MT%.����*�eӽ�};4<|n0�ъ.n?�GI1������s,$�E���:�9p/�1�3�O�|��VJ.P��ٕ�h_�:�<�Č�P�ń�T��b���V�O�w��6>�l�k{�2���d��=�Ŀ�v� ��H9J��O/oqc�TЗi��.�3i�\Kw���dmw�js{��w���>���r��a�w��9w��=�m*ߛ�(`���a���}�����/�#"]~��?n��2�US��xibr��6]��1X'�Ap�'�Q�<��i>�,n=���\������O���z����F�;�s�s�3|4I4��W��OV����g���uoJj���vL���~eKG_h�i�eT��d~N��ʞ�{V��1D(���6��5y�O4%zU��ߵ-eB�w�E�7he�l�@5<MVȝ%{b�J)��xF0���AA"^�G����Ȧ����������ꚡOV�wk��I#ذ%cRg�/l`��O������WBJ�_6IG�߃�v�&���3H�9�� �<��6��^�8�8[_�y���z��@�y�OYwNڈ� ����V���'�K2P�+Ln����n����I����x���i>������|�
�w��Q��տI�e�Z��x<{,~P��n󆌉�Eڤ�A3)��c��K6��s,�)��I;J-�gHĢ9��I�`6�gTm7'	`���Ї��������~��<�zby\������s,�*H9[oK[0p?���0��� �GD������Բ�@�Gl��7��
�z.�1���>(��͘B�.�(Kw�LNi��G����:)0 ����ǒQ�����L��fS�'��sD�.�O�KC���\qʷN�h_��\�Ң�Z��	��;���Sn��S�]W\���w�@T��(/33)�d��LV�6�'x�n��A6f�<���$UR����nxV
���a���By	L^���+M�\ۃ3��x ���� ZY��v��Co�I��p������i�x�1ca2=#U!��(ϛ��8��>�O���9�C�?����[��_�b_.?��U�0\��s O�9�]A����I�x}IZ<�'�F���+-u���ͳ@��.�(���*^@/≠�󒙛+ێ��ä��"2�͇����[$�1N�v�2�U$�1�k��jG ��@bGJ[��]*���S|�>?��?�� ����	�<�����/���D��=���?���r�h�x(r}�{
w
/��c����9�u�	rѮ��Yt�v�a{5��,"�*�_*����s-�_��QZ'�%�Ɔ*�sZn	T�=�����;8ޭ��ԅo�W�����]�&��f۬��<+��7��w�Ǐ�ܼPd��#�:N���;�`fժsB8B�c�'��u��Y"�!&qIG	2*s,%��%a�y��Vv�1���v��\`.���}:���2���adϴ}ӳ�R�����h��i(Of)��V
A�*�fO��Tf�Qg��I�xy�,�š�+���&���������^�M��>ئ�t�{�/qL9�t,��ZH���>N��3Z��ز&����e���db���h{�%�����*��ͤ��5?ǣ�����"���n8���Bݮ4��%4Z"���os��9��"$���J��JT��3P{�nMI�Ϭ�͑�CX*Y�ӂ���Ն%�4�#a�)����/���q��1��##^�7�Y��zuK��$�ʬ�i��������YW4v��L�ȓ���/��\{P�㟑B�ޟ���w����S~�&�Y��ûz��Ug��w1�I�พ�⯼����u�p��w΋?Ϸ@_��R�=����	ś�ݩA���b�D@����RM�yԀ�D�Ϥ��7^�Q)���	��&Z�;XRSzd+ę��>~2���{��[딮)��SE��R�ݥ7͜��R��hn���J_<;S2I�������Ec
3a��R��x�������y*�8ߓX%�%li
J��Q=}mj��]ذ�,��=�S$���ѝ����A�Vj�8�5qY/<{�U������K�H�����.ꙮ�H�'��{bPX��0/��S���bHp稲S����tu�@aL�BD�]�r�t��Ȩ���iJo!�����-?Me�0\tp����U�Y�+��0"��<2#,كH��>�������}�6�}�"\���
�ҿ�E��E��t����w������C�-�~nF����k ���P_���}w�v-c���y�5	�~�Lꍈ�v������1�n}�����"{4<\�+��<�z�����&��<%�?���a[�
-����&�>��e��[�s��Ňp�#���Y>й�@7]�՝�1��ff�v�L�e�n42�BȀ�`�D�v���9��@�d��%[(�f�d��OZ_�E�}£�V�"��}��J\��M�䧵?���$��l�腡xk h:˫���|r �=���6�*�`�b�l�++-	��wg �5�U�~m�˸^���.Fzz���=�ap��r/������j�{0�� ��ar�j,�s�ٗ���V�Ǜ�=y��f��y��y�ͳ1�C��0�-i\�]�|#���DZ&�NfyX6)Zp#w���!Z�`��]�ّa� ��ߏ��8*fԊ���3��=iU|��K��K�«g�Ȏ;VV��ݿ���æ�Q��(�k	�Ok���i��\�6��{8�wi%[�{��iۣ�%^�i?sƂ��^� ����Z�ϭ��yDI�ʥ"�I���+�
����8�0�0,K,y��#��҈X���ڨ�j����'Ol������;PP��y^���܎n�ç�L=D�#O{{�ZLcf�<���ܘ8`L~��J�zWǖA��SwOZQU:f��9w����c���w��^1iUS'2��5��w@/�� �*>KR�4�[M���l�j��W����J���p�g$�ԛ�Ύ�=�oK��.|c�5�_~XY�}h@IbR	1Y* H|:͌X|�P:9~�Y?Bi�5�:��"�b�Z�3(�a����ҳ��j-c���%4s��V��H6�g;il7i��I��5+^$G�GH�(vu}��v��<�i�[��^_�Y��:�'��@h=��'+F���Q�RWT W�nLJ�BOp�WTU�O�9��,�[�4� U`ퟨ����~�o<4
R,3F?�O��Z� v����dT^�z=-���yhK���Qe
��Q�2~(�$�C������8F�MҦ#&}L�b��3u��r%���4>/�/�A��(q3[)8`4�6�y�5| �?�9�C��h8w��\���?�γ�ք�Y�]�,nQ�; ��8���t(O4��*��xGX��k�'���2����~�=�Eݢ��h�$N��u�M��!I��Wl6���%�&�_o�p���I����l~�_�+`�jt��q�Rn���h�b��y��:B߻���Z/�Zh���cTC`�2ٻ;�RK�Q��*�Ld;�9�)�!�!�hS2&�2ܮ?��/�{�\w~1h��c2u�F��*��SQA��,��ل�j,�9Ա�>㬺E'i�(�3�5k���+�"�΍����|��#���ן���E�{����o������"����J)��^~Y���Mqc�,��*�kt`�_[\�g8�g���S�����WA�t�eP�=<Qoò���p�+Gqnx��mOq��.Zv�גiSԌ,4 �un�xyb�,s�(Vʑ��)����!�E܎���2Ԗ /	��w��*�w������ϲ�~t�Ks:M�b���׷w��	�H��o�af���2��#������y7r(��u:�1��練6LM��nx�FIS&f�O{���UF��le���_��T�[{��f�����VJ���D�r��~�s��<�0� УM<5��s!�Ŝ\A�o�W�4)O�0���>Ȉ3 e;��d�i��SuqKO�'�	ʙ�<M�����h�l�-]򗥟�-D�吕SAP,Y3�k��;�L�X�Z/1J'W(��-�p������:�HD�����؅F��s��vk9�$	.���8�����y&n{o�Nן���(�=��HR�c�5�� xBT�?�َ�mϒo����5�î�0}�2��Q"�A$ރ1�-W�����J|���&��J�Q!�W�kC��y�0e�P�[ϛ[�YW|�)�f�U�)�L�|a���-���).?Ъ>Á������&��ò<~qz%�a1��<*���vx��G$�c
^ő���h���"]����0�J���l |=,���ޗFЦ��>Ah�Ɲ9d��]�a��f���g�z��)����6A���J=�(H��*�4þ��u~���7�OV�*>�f7�އ.�Y}�@�� iTQ�n�gQB� �hoL�w�H�NB�%EA�}�ZAr��=݅1������V�e�5��*�Sl~l����b�5bˆL�>���?�C@�4 ��������٫Y͓�ɮ**����?'�sĦ/��H��kt�.��\'�/������1c]���OT�4�HbS��0Z�{$���T�K��v5��K�Lj��q�2�{�z��̆�:�!�	���W�-�F�����WѺ=�˲]|VH�j��?ڟ:|v��C�[Y�;k&,��-�KLm�@B���+P͌l��`��ƍ 9���G�ƤLtA���%�R��4O�5N���):��� `b�0���j|�p#�{@["��O�,�g�h"`s`�����u�&�K�fl������Yl���n'.�#�XE����U���_�e�w�PF=�}�em3��@�}$)���,'��xg��[��Qٵ�3�"�X�V�nh��5�'�������Y΁f��M�,X>�$h�Q��z����mu�ԹR���7��t��9�Y�g�t�ِS֝�w ��jEN͹��⢢���h�H�x�G�{n��R2.h�LW�So�>�X���=��:7���5�]����!F#2�W��é��/�icx��N�;nE!T-�锽1���)=N�^tĘ��Զ�Hd/��S%�KT�7	��ۺ�#U�Wp1��9�o�N� L�#���+�A�4��x��fӯLi$�Q&7�t�@U����,��(��I�Y��:y[Яf�({��k�xZ�NİC�*#��KÆ"h�6�"a�呸���ܕX�&k]o�14���*��z\���5-tM8��w���u�b�ruyެ���=�)�Э�i���S����N��M�&jz�i��O���T	��}[�T�����]TkiM���l&UIM�3˒���=��Q{{�����3��եOQ�<���qob�"YV�[�6t��������T��֮�͗NO�W��87�܅�T�)����
�nA$�c���'�W��N���xCJ�`��4��;r4��3l��fgT6����.-����_:�����|-�����丛��6g�,��-�KN�3c�k��^涹i�V��$�%�����|B�-F.��u�=���C�q��X+�}���o6'zꨆ�Fn�n�vh?Pٚ�N���D^_���KDbP/pỗ�﫛��V�>���b-i��Y̹���{�ɭnZ!2	w��W9o�&�k42ug��37���7h��\�Go������\r�@�H�*G��OiΩh�jI�J���Y��<��R��*���[�(E ���JqqғxZ<��2�M?��i!�i���xk%=BK���!n�1bW��#�G��ޙ#�T+	c�m��q�jD��G�.ʟg���]b� $|*���eX�xRs�gHC5�F��7٥d+����nN`�"E'���s�F��H�����E�~_�!>em�et���x#��o�EO����{���g��i��pޖ�ܛ��Mȡ���X�O�0s%ACoU��uMĵ�,)b�INhKC�oY��T�9��7�b΀�b�� p��F� m&���#s���/:;5�:]�3�C��\ް5
�1z��Sx�9Q҃Ar3~Y0���9��-�.�H&��Y��w���tM�c��x�mCw��W��ן���<�Z����@2�fg����^a��n&�(��_^�����SU�L�kx�[�h�o�z
4Ԋ2eP�[-S���x"��--�1����P�+o�~���X�v�|���^�x� �0�\H69��c������`{�(��~�+�V�؀���&�<�� ��"������x�ݤ����hW:+��νOX�xy-R�E<�,˨da��vW���}�V�}��or�o͈jp�	;t6�t��W�H���u��YҒ8�gUZ.�q8������_X^��l��-@��+�E\,@1	�ͩB�u�\�36ExE�@�4Vea}���gx�d?B�ޟQ��ǒƫ�y|��}y"p�29z�w��^�-��Ԓ�I�(ꦠ�"�\�v�y�{S+��xQ�Q9����U���&p�Wf��R��.�q*���1aRr�5E��6�Lf4S�5a��5��˅P��-�hf��`	2��E��u���<�ym����[C�/���HC"���:����x��.����U������ 5m-�*r$*i�g��B<,���X�� Ej���.	+g_�ٜ��pmwF5l��V�D^�iOۀD&�;�T�w��D�a�4�Z���]Kw1����l0Lq�G�����X
�?]vƀ��_��u�9���' ss4�F�⾦�]�H�R�k?�}�m���_�,w�')}U��[����]���)���BP�_(sqr}��g23=�xr)��͜�k9�?+�H�W1l\�Q�F��_�V����!2��xH!��"�x���0A�����nA��^ӎ��RS�t��MJ�p[� �1N�����!�
h�[~p���cT�t��y�m�
4��~NOG�V[T|�0+�ѓ!��E\����w�s��@��u��������ԭ11{0-+�L2�2f�L��.\~��z��V�)�t����г�@%ާ�{��1d�f����f^����7^k�7P~Vy�>-G#@�0���'rlvX�ݚ����;��u��|(��n�އ�fxiֳ�d��sv��2��\N��礤kv$r"��;*��Y�9 &^v蠙��.����6�7	@���0��=��}���b��+���:��rr�S.[fI� �-	�H��f99kS�%��~��}&ْ���Z��՗�3I�Ta�f��L�g����N���N��a9��qJE��DIaf9�u�>=L�O�jL��e�j�Y�Hs��M^���؃pY��Ai���]��VYUg؈��/������ )3đ;�L�?��/�O٪��k&a�Dr0s��W�_C:V
�J�<o��&�)��Ւ��`��+���FA�w�_����H��͡d�e�\�̑W�
7Iܟ.��ār
��N�����(R~��g�z�T�bK�������~z�W�h�t�^#�_��V�t}Bs��I��9=�U���1 �2TX����í��h�n<��B�+���h�p*�}���r�0@6��M��̧�T���X�����c	��B+p�S�$����6����J�R.��L�~� ��;���o��D��٧�3�u+��_ցY�����E��+�߯0�����hv
���XLM/1?����[�W�)b�i�s���<P�W۽��78m��	+��w<�OM�^��3����;z��M2� ���s�3�AʇB�����D��_��{���]�Ծ�Zkh��U[i�5����Z��,�C�P������y6"5���L��LlU�љ�s�s}�����Gx�ɠ5{�ݡЩ_)��\F�$�GEƖ�J!�=T/�'���Yv��b��@��d��5�������1�0Ǐo����$!�� ���U&�j_͇S�-:�1��U�\�ј��>���򼿁�Վ�Ρ�8Hr����3�M��q�!����� �hNTdX}Cp����1q�~t~y�� Ϩ-t��V���Yu@+�*mC#:='�R�����#mfZ_N�z�b|*�'F�*�D/
�������6{�~Қ���{�~ ��������6��2w3�
m�M����;Y���ŗ*�"��*n ��F4k��v���^�h��x%�F�0ؠ�o(N��p^)+��R1!S%�}?���?��UX��;�JV��/{�e�~cv���Q
O^�p�E6�m/��#��N9`<F�/��{'��_�l�CN�.�*Z-r�;�?r�}� \pn�q���G~��3?9=
e�5�}���()���+Q�i�0��)4������O
p�/�N�:��0�)�� ��r��� �n�]�@�݃RbW���$zg'w����38���Y7��aʜ�(9iYԀ
��y�E��ii�����]�S�w �m�#��.��h��K��'V�6Mȗ26K�|������8b���:�w53j�зw�t�<�zteQ���xYuL��O�2�_ʭ?��,<c٭u/�7n�/�T*��\�#�`v����Q�����Sr�<i0\PE᪖�xt����Ӣ��:Rلt%�p������y��_�i�a��2�:tqD��^מφZ)��g�)�ʍ��c��&�ɋT��ϰ�k2
�S2B�q��w hS-�.p�wۤ��XxD:��بm	*8[^�n�For��)��8�e65:��g��*�Y�F�{�S�" sg�a�/7��s�+9S��і)tR�a';�:{nc�98N�K��V�`I�~�����'�B�Ժ����� 4��S^NA���X����g�paE��2Q4ט�{��{b�?<s��/����ͻ����fv��:���J��⒬$Ks���$4�C��ڭl�eTiz9�j��L,��ɴ�9��s��>����*2p��/�Sܝ��ѡ�4~���2�WGvd�˗=E�\���~���X*�$��,�ĕ�#�xG?��|gP�,�}PG�m��V�Ŀ,��Grp�a�D�u7����+�@�'�.\N���<�=Q||6}�hnH��$bzy���ЖԤDiz����)G�u��
x��1re�+����
����}T���w��`�ar�jq��K���ax����I#�Hp�k�;FE$��pw�R��p�m��xJ�ί�hٖ��m��q���<�+I4������U�}��O������Kbv����9orrI��$�\_kn+kAviW��ٺI2� M���?S���?��W,� ���('���0M96���_Q�TD�!�Mƃ��d�eO��~)M��anL�Mz��9&������!)d+�5+�4Ҵ�ڗe��	��� & ��(�5l���2���q4���Ƀe���¢Pϊ��#]Y>R�էC��ٶ"���}�ZEJ�`~.�@��B`���l%&���)�)��e�ȫ��ے��7�g��� İ����,�v�l����{����6�$�-9����صH�3�2O�mY�ȝ�S6oh~�ʶ<�)Up3;���;6��n��R��l�Λ�Љ�H�/k׿
��U��J f{����4�.�/bn��;4|lF�v����>�O]�=;�^�c�,���k�Ȝ�Q�,L�ba ×��{�2��WnTO��"Q��J���j�I�x[w��<`����O�$k��ѝ�sL^k����M��Hs-1�P�Df��E�&)E��dϕ���?Fdz��L�Ks�>N ���ϛg���a����g��21���{S�f�Aŷ� q�7������&'gsѽ�YS��m88�H��e����O2oh��*�YE8D�io��q�`��\7��%|�Ǯ]����Y!��Y4�D+]=���BخY��u��~9M.s���"����r��9S��%���a�%���(�K�[��m)_r�N`��ْ4`2궍K���c��?Y[��B��ٜ��oT���cd,�ĴT�.6�H]Ϙ�Q��	����XxS8�Ғ�nǠ�\q�A%	5� ��A�<�@eH�LAlJ^ܣ��Dޡ=�k��D��Y �:�� D
������?{G^%�hf�|3�wۯF����� �q��S�K�Lq6�Qҗ�yڌ/��ë�u��Y�Nhej�'s�[`p�P�@3�=�V��f딝��Slӓq�_�w7�^���I�'��̌"��3��C� Ij/�G`�fc�iɦ:�GF������k-�e�Гe���^�pk%Bv��V�����Ϳf�0�m�T��X��(wؙg+F��OVU�I���e�iǙ����+���{u��8(�qk���l5�
��6����/ɏ �Ui����v�4�&�����E�%!�9p��</
j}"U��8����c]+f^{���S���Բ�fu�W�dϛ@�E䕪L߻���m�s�M��7K]�[{��H���`�3�����S���m�2�
�\��ϱ���d�?�7<v�[���?}�ݭ���L���6=A��YM���&<|��p $Fl�Q��h�b\j&ZӞ����+�+�5�D�N~���Dw
?��z�w)�T���q�TH]!�p1��{B3�ה#�;�5n����w���]]�\%��;d�AR�x�1��[B?c�m͌`�p<�"�P;H �-�D]�j�*-/��@�U�YU�S^�UV_T�g���ln��s��\}���:]�<z����E;�DVd���#c�!X�G���(<WS�/�Aց4!�J��(F����֯�W�]�WU2�/KTfd=\�8>6�Cv�2�Q�+�h ����9��<�؅i����@WП�o�,�.y�a;��8\M�D9^��He)TI���`@�yuQ���Uʔ{@Y{ul��<����Ǚw����*]����p�ʎ���Ahx�b鶓�̘���ɓoM[�z���ѵm�7��C_��D�:��'�y˵��x����%pu����l ���[q}7_n.�d�B�+F�A��v�ap�{�����՗������k��ݚ�	D���7�C���"ka^`sc�-�����;3�^�m,/V/��M�<�<EGL��I���U�p���#���eO�,w��..�����E��ު������1�O���_�IƤ-��F���hv�Z己�Nt���,v���Q��e�=jDΓg"*H�,7�D��2������Qd��d�,��nf��@drB[E��ן�i�Y]L���ج�S��xR�&�-�_��Sɢ��쳥Y��"%IkF���<�3���ol�m��E���He�z�xB�`�sd�� n����nT؜�Ǯ���zqV��`ʷ�go�4	ak?K�/k��^kɚ�W���C�v���kt����Wcs=���p��a����$�[2��49�
1qm�V��
���TO;��Y
����oL��%:D1"���x~����q)V�&���+Zꈟ�W�u�?��_��N��H�~@܅�/톩�`Ӆ�q@d�$be� 4+�	�������g��U��U�ȧ����;P�	�b��܆!G��)����X�H]�II��x隅S#�^�c�%f��t*�WVCQ�4���f�=��_�9� �(�w�L~�}J)e��b��Չ�!
�% ��Bi���S�jzyegN��y:l-��E��&��L�f��!7�k R���\���Jh����)��$��g(��iQކ�#�Q 	
��vry���C���9<|�)D�i��g/(��H�B"CTZ�`EY�`�eȳ!�l�{���5+���GL9r�.43�-��ʹ���p�D�B��s�a}d���Ō����?l�mL��,�\�����ߟ��e�nf��x[��p����C��&���U���lT�z+���]|�����ʞ�%�#)M����+�BkxX�.�Ğ���o;z:f)��j������)����/E^�o��y_@�G"]����m:Jy��1���#�����S%�m���� ��㛦.���������.��&3{�Lfc�z?����n�u���r���m�<�d�dd��^G��Q��%]�fe����,w�gg��)���Sbû}7
��Q�	�*8�n�:�
Q�c���E�Z�M�)�jgLko�v���g�'4�Db��{���+;�4~���,,����m�i�t��1�{R����mZ�F>Nj�թ}i����w�&
,��W���� I�Ȍ���!��U�J
�F���e��C����W˒���"X>*n���B��`v�d��a$��n|��q�+�Z!$p}/� ���]N���8Y�	���7b,?vS_:����xo�a/䶹����ToXD�h8��ؖ��'|=4S��*���yܤOs/�d�'�M��@J��s �?����Od�UET�Z�3k�bx��HI�
 �,��Vw�"i��
�Т�xs���:�ƈi!��)�3�1�Oq� Kʗ�M������ŹE��Q�����R�@��E]�?�f_YL��8eK�-��g΁^.NA�w����r�G ���V1���Aø�ޢO�BB'�o��Hr=l>u��q6��*�-�ߩV5��6�/L���\�S�y�u�~�k�O�D����*H�T�`�4{+�O�G����+tP9�ݷ���Kd,׬�|c�ʠG�w ������䋢�˫fbi��X�k4-��1w��l������Ek�*�JbԮ-��{k��GP�(�FĬ�gk��"6EQ�h�h���+>�_��<�s��\��y��>׸#��Vh6أ΁`���C�ŏ��u��������*�f�+�&"a�i�u��� �1b���$>�^�cCW�D"�}�N���泙��]��>ώq�8^y/*�drZ>�n�$�����'�:�":����%&s�,ڸ��J�F�d'����s��j��z���TS}������186L����<��g�c��dl@��8����(a�DS�������ӱ��c_|q�c���Ӝ��9K��e5�,_��F�tl��4��Q��)5	�VY��hG���b*�X�M�Kg_�w�+�{�M)��[��/L�)n�s�1�/Ѿꕪ�����Gu�ξ`���լ�y|A�ӿv�C;W�!����x[�?^L��./(lG�����a��Ud�։28��^O=\83n�am/h`"�W16��B'����BN*���R�ot��-��g�P�����hI� ������6}#�g����� �(�:vxY+[�[����.�Pc4XV�iA��f���/Mw�lz�H��m�j���&�-%�J/��]�/�M�c���/1��y��?$xMr�.� �5�1�H_�Z��O�70\G��	)l�<�;d'M����4����X����ڰvlw�j��L�;#���m`�v�jr����;2�;J����=�#g��f�w|���~�Z�>>ف� ��G5����A ��Ppo�!���VH�M�ZM
��g�d��6��z�� ��vV�oʝ�KrQd|�s��F��:$x�ɕ���](Ьm-{��2G�'H(�퓁�I���k�.�4�Q�Ї�3b ��cVk�����\��Q2��5�䖋)�鉋�c#�_�4�{?B��lԚ=�)����[T��c�l�IX=ǒA�:�Ch�ؐكI���/d�ߕ�G՟-�n��;��F�kV(|1��M���H���4!�I�O#�5�w���QƻM�����*=kfz܈�ō�sW%�p�gwߧO�Q��(�����M�ԫ��,��m�-�C� }�z�lm=�a�����vO�{22$k����a�G#,=ȸ�`-þIl}���³C_w���H����M3�]nC�v���V�Ef���jv��{�?���pG>��*bW�h�j�����;��}�/� ��r�EiYA�剫�6��I�hUM�ڂ���k~���.,�U������h�S��Sb��̬���G� ~��T.u������7���u�|��)���/~�&�L2sBF�V�Y;w�s�G%���<=�n�O��ǒ
}�d�{,������gnc�"ji�����*��Eg���Lx����TY%�J��&����P]P�j�'��͹�|(я����Ja.`lW���H}���3�����A����N!:�/t#$��5LD��#5	t�*]��ɏ½�]�kE�o��T���kJ�iD�`�x�fѩc,6��pH�ګ��U����%I�&HJ+�{0;M>~V����G�U�ޗ�������i�OفF��=J�9HS$/$�\�'1��{<�A�K%+2R���ڮ����f��;[<;�?��O~�e�u��nF�n���.����2�&�Z$+�>َ��}�9 ��^��j12 �ޑ���'��0�3r���u���α
�SU�{�m��;��W�V�b� ~?c`p��|�3"��d�_��A̗\^-jgkEѨ���/���&+���ܷ�v�xWO���n�ɪo[<�w��w��ӂ����b�r��MR� ���K�D�����d&�!�鵭%��ql��=����j�׃xiImE�U��̩l�塯��'Y�J|1N	!.�EN�k���:'�F�8�3O�C}%B��)���ӽ�x�\��Aw^����/Mpѻ�?�$��	Fs���Ս:�[���.G�{.)��?��{��f�~��D��&�'��e��G�%�!g��o3�X3��>��b��n������f���	k�8�K�1IӃ>�-[�AD���܌�860ʩҶ�JО<�_i�[.Oz�2N&�Q��'���:�E=ݝM6����
U��H��
�Q���˫<|s�Z�L�EF��dN����3�c�R45�^&�k�qi �6<��Ek�¶��XA��n>�}�����x�b.h���T�F�� ���pQd���IDw\���桘}d�k얹���3�TQ���8�չ����t�?fs�;���=����+���LaC,ɷe����&n?�sRJ�F�r�i�����k�=���Y�`���e�-@(��b������I�y9u硬�7H�,~�݀LZ r8��1�CδQ���x[w��)%��N�{�be�g]��\��A[�/C�ϙ��o_��x�^]���}� 3��?���Bgc����\���st�����
��j:�ߓ���6y��Z�o���-�H!�$��}�����|���F"/	��1O��i�� spǳ'��B�[��>=T�H�zS5	��$���E�^ֺ˫I����V��<c�R����ES��Dm,�i�I����w�8}~ȣ������:N(0T������N�M�!R��=�s���n��mpvȻ�9�.�X	Tt���^-*%�Z��߆� +���b�l�#�_����Y�|� �9��YZ"�'~60����3M���/���1w��H.w���4�����^���|�ŘV�1��o�/�O�+�3?P��a��xT3s�
�}w��â[�+[�'N�ǚ1�Tw�zpƃ�y��(�?�;�q��`�>h�-�;���<H�4_�0��I{v��H�lC=9�HJ8�S��q�"�D6�5JƠ䍷���3������k�|W�E��N�B���p9N|�	���x�s��B]��giBUz�vܸ�����nC޾��>)Cn���u��4�<0����Y��Gkf&���W>�c�N	#�D��sY}9;�nHfT�sH�]*�ʢn�,U������@���E��s����x1"D)|`:<C���Ӏ��`B����2@w��8o��s�����	IT�?��0�/+���j �k��s ��}i<��ή�����G_ɹו_%�1�:y�g�H��d@zS}ǎ���;?{ea�A����m ��K9e�6�\dj>d�H��óf�y~<�Ji~.��b{U`��$�k�9צy�������k�& �������D����Zw��y:aƃ1��PA{2��q<�����unljG6�4�&9��*��+��p�]�aư{�.�TX�W����	�@�<���BT�Wv6�x�o]�ٕ�آ����~���('�������ye����습�h�e���s�ӑ\o�d����6{c��cf!�n3C2��@�ɕ�Q?sS?�L39�j��0%�fh^��ܽ:�����͵��ɜ��}7�B	��jޞ��������l�ʔJCU�2��\�ǆT�ǖ��L\����?c/�t�{,W�v)����xJ�7H�^���]˄)ƺ䜺��"���@s��m�+8�yz�t8�8�hY�!�7V�V��t*�fR��ER��M2��n*� �峫0�ք�ɍ��DN���N����E�Ϋ��Cئ(Ѷ�sAH'�$��+�oM��k�>Hk��A��$�jI�?��CI-RB�f_ؑeH�Dgj�ȸ���^�yky�Yz>-\m9�0j�K���U;<�rQ��Q��8e�PЮ�-Q^Ӊ{*Q1Xe���K���h���@}UUw=�?���FM��B�8Ѿ9��G�<o
��,�H�ѣs�����SZ��f��V�|�k�j�U?ݖL�?CÄBZf��?�xv{���Es�~ U���aڂ�@8q}e(E�;��t`�et>����r�M	�Y
b��e�H�j���r���o]ߩ�1����w��x/o�pbMr�&y�Y���J|��5ޅk�ܝ���t�Δ$>�0��<�T7C|(���J�()�+-"]nPh"�1��t�������V��>6=w|��3�>&���wSf���+Y�Yg(N'��K��Kq<�����j0	�p���^��\��ǯ��&���qd��n���.fn[ݧ�E��A����\�q4E[.��"� j��o�m+�K(�i9�"q�p��&$K���݊��3o:^⬥�-�UR���6�+�s��#��+�d�yP�- q�� ����A�F qu�[U���wc<��`��������֩Fz��;Z��-ܽ���K�YR, �~㯟�z��9���p�/�7�, H���WP{u�2�j���,i��jA��@-���Z�����E�����+}m[��ѷ�2�)6��xd�h��3��J"�t�<�Y�- ����dO�iNO�I�Hb'R����[���|�ԅ]�,����%�\��RȭZ*��]"rx�{����<�L��Ӝ��[~zQK��.�9�g��O H�t_Ծt-l��]}�.��9[����D��?�;�k�H9�`uw��LcثJ���=��	����q3p�.6������<����̚�Dې0b���s�}�]�Z���X\��|�h��ǈ��fȒ���R*ǿ�|���[
)x7w@�$���yf�Avm.E��fuJ_�Ƈ| �����j�G�>=g��"?��������:�mۤ$2ym(�xD����q�E����h(�=w�h�Z�s�곌����<F�h4~Y�[;q���)&�u������tZ���GH���$0p^��3)��d��Bm��.t�,Qܾ����/7��6l�P��3X`�����C��d^����� �9f@�����~�~<�x=M�k�i��#������r�W}$a���iė)�|��#�Q=4��f	I�����i;1E���zHM����j�v	�ܠz�W�G�12�.rL��]�������s:Nx��vDZ�|(�*�j�	[�"o2��<�j�n�N�Nk6lu=�$<��K�zdwW��XH�Z������L�/S����/���8]�E�7ǆ^�,��c	k����G�[���OyBA��7�IX���7�H�S�~�`����gi�B�A�)!@;Wr�=�,�{z�.JLJ`���{��4�;a�R={ �DjU^�V�������X�߯=AlbC�ާϜ��?#�M/�u�M[�?9�����C�  |��l�D8(Gz� s�bUӚ���H�x��k�����I�'l�8�ʵ�*��h�=/������o��U�Ƅ[	��`sA0��|��}S6<j� hצ�����جQ���x��E��Pه�z�����婓�yV0�Z��+�G��;���[�l	�z��<У��:�6��gTP��2s�"��Mk�9@<�vI;`g�(Ȝ����ǟ�|�U����5��z�w-=-�
�Ut���K/73d�䚭�wo�:L�ݚd9o�~��M~�����տf���t�}�!���mيk�Yh�	iJ�-"�:_M^�x�%�~�s��C6���or@�VW$��� I��Q��g.>�St����!��,ݼ4���yO�~�?����,eX�4��seWzr��E����|�[��v��)Y�������]��w]1j�<'>�Z����e}�`�D�>�����A ^�f9	W1�lFF���x�-s�Z4{Uph�������{S��C��"|َ�T!T���:H����w}偬=�L�L��M�`��sϐ�ɚ|��Z��#yB�)ߍ��\���:�X�z{z��gC�ٗ�O��^����0�0ܔ�o&rF!3�5����[6��πȧ����M��볒��E>�w�N`��6�oP!K3{���T �[����o��@���(�Jib�٧S����y�!�����E<��{��$���Rd���Z��Z��#,�|�S;��R6	&v��c���fqg�A^�U[���n_�����*�Xشʔ�w�����У�-s5�f�5��i��2�7����E�]�k��74M�#A�������@�_�|�צ�˗a�x�66����꧜<���2.�	?*y9��'�jR
����8�g��D�W{V����J��i��^y^)^:�E�,,G2o$����)#e��>�k[����^^�w\
��.:q��0�{��9{5���eg���~��f���v7+��K���G ���S�;���9k���5T���{�W;��*ڵ���Ӳƚ���)UK��/�e���Y�4�iG�4�ǁho�QQk>;h�\��l��{�i�$�lѠ�Ɖi�������,��HRN��a�:t�aU��|ӕ\����[y*��`�u��u���~^|M����+uK�U��æ�kP���y���^�*� �����vL6�XI�����|��M�z���u�,�d���N�CƯ�~�>�����u'���'O����	�R��0.�h.�tL�e��".>���(d�����
����\.�rPBa����W��P�h�^NH#�E1R(��2w�����͡X_)�2\������#�����e�Z	�Kܷ\�o��I���>���Z^�O�U��;�eQ���H�� ��z�r-7�s7��R�*�>�� �7OA[w]��Y����i�y����y���l3k�^3�����CDl�BQ���/<�樨oi�����)q�gA�R�<���!�qj�bLr���g���7
��V
jP]��b��Y�\s��(ޱ�o\��o�d�D����&M� �m�8�?i��!ݭ�� �w5_���opq�_]4^*~�<��Y�Ŀh"ވ;~�`Q�8�OGi6��M�����vҗ3s0,oHD�i6T4w~���ˉN����(�|�s~X)� ����*wȅv���o��(ؑ`�4F`M�0\pZƥ�fy���Ui72�i��f\�S�	�9{^A�|�FY�)��m� E<�)��a�������*�O'�U7&(=EP&Mju��q�<@�/�)�{���߃Y�}�V��Z�B�������É��2�Z���ǋg��8��
�@G��!���yl�}�/36xW_�Տ����)^��R�i�{�R��j'��<�4��v���G˦�]E��?0!�|��۳�K�|X|��@A�W�;O�e�N_q�o��:siA+�;�t��В����IHs��q��$2��6���Q��D�RFs�ULc�@���h��#�!�C�Y�s�.�lC�TYH�ߜn-V���˨	u���.�|�Wa�b͗�R4x�By)*�)s��Ό���M�4l�S�����tsZ�UE�s��r�����<,�&��L�DYLk�N`H���&�9�b�^������W}#���Z����� ը%�0����;^H7?t',8oTo���������$w\I�?o�-��"��(�wЗ*��`�l�y��	���p����*ɟ[��R�>�j:�����B�[��{�v����m����i����a{�Qz1�9��6(�4N��j��)C&�Ժ^�R� 0��
7�z-lG���P�]���;�V�7�\B���F����Q��)�o��;f�-ⱬ�6�v<T��Ҫ�ة�D��u6�s�^��!�9�������P��2��2�d\�$ha{�@�#�5.*g-!wJ��g�E��*{�6��;�/�Q������$��=��%�"lNI��u�O��D�W�- VeQ{�E�Ka�v�y#���v����"��e���P#�\2��g���r�W��|&eȍ.7�Z����۽������t�u.ը�R$�ML/NT|2R�|'�q_[N�鐦���2���bB!8�	��}a3�H���,�w��ʛ�X��t{d
~'���? ��w���dԤ�<���pb�I��}"��͞ !�?�Ͷ/ʔu�`A�_�SM�d��e�e��j$�����>YH�Ҋ➺\��s%G.��MHa����M�@�D&�E,�&�9�,:�zA"�&��&�&��#i��x�_�`��],"����΢��j�E������Y�?�w��>G�w���5��N����]�{kq�u�����j��.,�{m����K=hh�sm�#�x�2�w��oU�3W���i�(�q��������I��a�@�ۃ��c�����Pz�pG���aqǏ�-���FeS%x�b�?�<N�=Oq�k�5���3c�~�g�P,9�6T@�Ǖ�j�X[��Ь�p�Ō��XU�!�+j�t��[R´\�*�i���̸8h3��gZ����f?�ݹ���G�ϟk��l^��{��8�`�4��r�wy,+R�tT�J-ᅇ�P^`���W�o��/$f�P�e���|U�����vbF�@?%�C?_;��pU�e�E�=[����aZE4�v`Y��J�E����*"��5�d��.=)���?Q�'���xًM�8c�g)����^���]%�S
��7kي2˭&����[��ƧF����n��'W����8َp^k��>�W2�5:�@��M����9mV.�?c�<�pc�f�����kS��-�T�c�8�[ ���sp�ٱ$��[@"28�ʞ�:O$*isUo&�W7pw��"uܕ
Ԧ�O�� �����B�Ϻ�y���X���E���ݎT=m-.��6�����Ja%�8�|���ƞd�0ǔ��)u��_gP�����s���9ިT>�̗�$gQ��_
����i�&�^^�;��>x��|��G�IB�}�G�Yo:�`l�q����넡ALM��
l��lf��|�EqbI�W6�vh*����@;(�����NV����`q��ã�����K�m�]�������᱁�rp�{�"GYv�����P���&�OJ�C&�p[�Z���i>C)�W��:��pߵ��@��U��,�XUR`it��,� �#��;��&s���N��j���Mק�o�Ы����W��ũ�kW������6]�SCTh�eԴ�9_dm��)2!Ϳ�cG�7��C���[g��
a_pWߖ���V�;-����TӳkH��Om�T�ƛS��"��Ts��N%�~(;�y^%�;�P�b$�x|�8�uT��t`@vG^l���ٵn꣸���8�o� e�Vj�-�����3��Uh�9#+�M�X�Q��@���Nr߷�$��<\a��L���S#�d���Ы� ���2�ޮJ�h�o�m�\b ���K��ԝ����{�w\M}�"	����eG�D{(+���췂2��8��%�{�+�[���[���_���P��f��FA~}��p!�"��lϪ���O��X� ���Se��)ϩ�RjED�b�C�����F}�W��B�:��
2�|��j�/�w��ygq�@>�(.Z�B����<$Opٱ�xg����	�����F]�2���:w!�E��#�ZIu,�u+ V*�����X�� �2#�5�sI�|�/V���QHi�GسI&J�C�fy�}O99m{��bnC�e���w�3&�W�C)aQk��p	]�]���L�18�(*��p$��ԧ��*hb#��Y�Q �;q�d-m�.	�t�&ñO\^�9q]���r5������_�������Y5u�w�q��RSD2x,8��mȷ{Bl����mj��v��]��tso4g䏥��W��NM�y�H��;�^K��oj�u��'�3n>.�K���n�G��I�'�ĖF�/�����g-�Mt9Y�Φw�Ƀ?[��[�`ǅ"I2y:��$e/�x��L	ɡ(��ҨX�(�������r���I	��>SK�Wh���E;�r�ǡ�"ၒ��o�5\�Tɂ��4(�@��QYy��b��eЈ���}Ӆ��&my��.�s�lle�
W���f�/�pu���꒔\�Y���+J�4�<#E��UP���O�+�T��>��Bg��(!���j�\>�~B���*]<_)���[�\M�K}��P9^��@�t{�!&�Sq���T�����:oĻ,g��@��%tOt����	_�����4���!����[K�n7%�Q�x]��` DH<i�Y�٥�HM�;�	)���F2T!H�DI���ə��Z�R��4۟Î���e�)��jy�Xqy T����)�|�Jq@���0�&��U*�J�'>������#�t�Ų����&���a��/��[ �[.{�:�\:]K�	�6]O[���#�X!�I�<v&�!ް4�99S���
�b̎�G����<��
�==���f�9L-��N�/v��܁��)�j�^�9�.�̵���CQ�^f�1\� ¸wp��(�3|�}���a��7>�V��5iI��c�o(�캣��h���0jڳ>љ�0R��Eb����#_XT������'�T��®>ʫp2~���M�k(�U�<*k�L��ό�SL	���r>���x���4fH+ջ<���1V`\�nz�u�3c'p�~p�r]Er�/�t�.7�D��޶�C2wL��w�ŝQK� ��<z��00N���U�d2#���*(#o�?�	��j�qL�E�S���{���&��;�/��R���@}��� �V�o�kQK�a
)}0C�;��
�V:��w�_�y�J�H�I�Ȳ�rFc#�\8��c��+�X�g߷�611�:��q���irʇ(x�D���(A6q���� U��]�	q��[�	�p�w����(��	�u��Ϝ�����Lۇ�#S����Y���\0�^�4���*�t,�ߥѦV炴��T�� ��yi�!�Waal�UoX�O�0��.(>���\F�5b.k������;9�C����ܻ3�e�!(�=N�!"�C���z;����ɿ�)ɨ�v�A.ݞWr(��^Su��Mv���Ϸ�^�K"SκX��8(K�j�=����Y�Ln̩ؗ�z��*'�W{i!��S�8�>��h�⑗��nΏ�hk��Te��`��!��Ď�p�`�����T��S��Q���w�Y�<4��'���r_�?>:��M0�X�^i	}����a&������ti\��xm��I��,Q�l��贓���@�"���aMc�>9؛�v�n9��c2�j���&BZr!i-_}(4e2ir�L��}�9��#}c��)�W�.�#�gE����[C#�^���j>���Ŵ��b"i����� c(�Z��������(y'�m�_T"3���&�yi4V��sGR�0#D��A�+��ոi9(���9����wt����>�����!�3 �G�`�?8N���L�����v�Z�d(���ՀF��/�l���V
h
�ۄ�����DEȘ�����5�ÔB��7�<y���v*�D}.�"�q��q(�K����K����b޼'�x�>�(�W���f�3�k�G ?o��:�_�qps����M\٤w��{4�C���uw���6H��ۋżL!�4_�a�ǔ=�#��xC<���X��"K�ݭ��%��(���v���=����~U�>�.���Ԧ�P���Ϸ�"J�j�ڙl�f4>&;������~�^��~�qhZ|��P�h�g�B<���\o���-}Թu=����Ç��3�0-�X�I0���@�L0"A��� ����DWe��������x�E��5����0z��QY	o�ё�F�:��Ux���[@-�_����!=Oih0��'�J���~m��8[�����f���@����&2A�pl'F&l��1 �cM�d�[A0Ap�e����u���jn��}~�w��*��QP�'��Љfla܉$�(�&S��O_����VV�:����8�$��?�?:zv�HD�n���2�޿'�xw�%��`
?�kj��:��X�r�Җ7nV�w�t�MY�.4�� �ARsg��"c�I���p	�|���f���F��#z�����''깠����ç�����&�����E� �o�0��珆Ϟ�E ��Xcw�}�����q��I�KqL�Gy����h�e�Yɔ�w�����K\���a ����	��/g�H���C�v"dO\H��~�!c��d~wބ|\���jk
O4$s	�������G�^�+R�7(r�H�B�	��&�O�g�T7�x�����&��bm�w��W�*�PIO�et�/ot)��r��}����V�tI��Ɔ!G<w����Ś�Q<�\��EH�Ąk���x)��%�cK�d�\�F��\:J7b|�*�k��[A��f��)����ȩrc y�%���pt	����܍������T �̷�?A{f�T�і�<ۇ�?V߀�rD�����I����sn�`���&��3� ə7>��P鯸���{���"����K�V����8~,��+�f��� �c�sf��K�-��~A�?50<c|%�0���_�h���d�>���[��W�n�����vC�Vȑ3����ܣX,��@ 6��}�%O�&���z{��v�����qr��:�")�ל�-�?�XMc�l1��;mA���QWa%B9��cuO>��JdA����ɶ��a����8,����@��v,�?f���Z�wM�nX�p����������K�A+�Py'��������O�����E�ejK�	�q�O+]|�A��b�@�{�x�AVu�s�HT䋔"w��I�E��T��R$�{���\�����?G��R���AJF˔	�]���M�0=FSv��XTw��������X�v��7R��+uVΦ�EV2���w��?V����\q�I��v��sr0��9=?z��>�����b/s���J�sUG�	L\['�Y34�wZ/�8����$6�F�Z�)�]2L������R����M�_����ȈW��y�)�|�ׯ��f�`E{��y|�D=o�G����;m�ZY�O��oS�\G�]��6�����"�FkG�B�4E�m]U1���'wV/��Q<'�o��&�ktp' k!�m���f��胐U@l�㍭�D���So�r
@���h�tz�f�-�;'4����E*0�ѐ��w��T�	��
����)������3�X`����,��θ�r�f�)>MF��L�M�)��}��I(�� 33(6 &�Voc��bdd8�:��6�������г����{+>6x���,�[���6��k��7���iLT$WS=~4ҡ�z
4W���u�5)�>__!�΃�|- ���#��X�����T�L��k����5#a���p�����kl��>�d5�G���d�^�M,;#�88Ν�u�S
\�Ů#!�;h(`<(kUWh�'���`�j��1RTBvMw�?˾�1 n����[�9VID'H(�Ч�=V��3�so��cڏ�3:_�t^o'�_f�ÍD��E#��JB<�H��:U��'��IC�V:�C�W.��V~J�%$���|W���T��.���>h�8��*jZ�?s�Nئ���ת��.N���2��)���MR�����"��2=��o��T�O�\����2�Vd�p��y6�W�㳞3�/�&@�1"]�zA���x��_4��r2*��Y�
1z$�f�ݷ�,I��
���wv���'�v��C�M9���W i�u�B����G��/�Z��{��	V%0Z��@ox��>��� ?c�X��ƙ�ތ�%9�9�����m.��K���	J�瀿?�!"���	h��2��$b��RjjC��f����Gj޻�T4�J6QyB�5��@���Q_G���+�t��r$7�|Dt��|���������+�K9�z�L�[��ggW��`�)���PFN��`&�VR�����$��z�D�N����S�e�=���ȓ��h���q�Ң�hI�	�U��<��.��s��X�9�K;��!_;�F�Bnz���ET�2�T7F��U;ཱི�.Z]y�
�`
��ۀim�p��b�*D_�J�����~�Ù�k"ޙ;�cǷ���"O��|i�jQv�ĉ2Ն�`��נC�O�Ի�(6�����]	��yd���!W7���T'Rtǣ��� 4˅�k��tζ?�o Nh\��"�|�N���.�����'>__:fB��v,l�}��MlrQ�:�Wԁ����k�CBo�P~c%W�hoT�6)��5At���O?�g��}�;�<�B��]�Hz�n��$s?S�	°�^�G���vG!s�(�dSrm?S=�>��8����o�֨H������A_�|'&��مB_�	VɏP��_4J��f�my2P���n3������T+Hq�C#��������\����t�f���jWXMA>�<�i��6\��B���G��7�%�a�.�GU���2\�4��H��ųQ&a�+����⷟ɘ|׹�yap����!�"n�&W�i����"BH�G��&�[F�P��x}�K�vج�w���^�j�_�`/}�N���S�-s�GE%�|d	};8�#�3�M�4q6r�0|�U�3#����<����tP�fq�m�h1��m�((�"�\��.Z��Y2���A>6F�b��Xq-)-7+*��25�Լ��`rp�p�7Ƚ)j��H/���U?LXW��M����<�@��C�4o��p�𻸪Ud�m�n�̛n�t�4W��R�ʟaB�~&d(��jvֺ2�W�Z=�@'5sG�\��=��[��W��Ƭ���fo�o3s˥,J@5�D�Ɔ�q5�6�"���\{c{�NK�`&���������0����� �9	����� #��>����X��I�.x=t������ F#�rN�.]�F��uz{�7u�a����gKj�
^�>��$�]�53���_7�2n���5��Y�)��	���g��WS&۳8�09e_	� 9���j.=��2��_�X=��`��q�$�J�H�;vݽ��/nG@��W���Z�S��g�<�Qh�h0l~p�b>4��'��ڝ�euF}��<$�� β�C��S}{R�(^�]o�.�����m����x�9%T.��]z`Λ �S�ϜBڛ{~	p'�Xtм^��p�H�=[n���s�Њ%�-
4��r7��-H-�~\ܜ]�Ck	���9�����FF���W�{���U[����*��8�`T��:k[��u��<��snB���Kt�=l��m\#�\|R{��oOM��t�6����Z=�N��ʂ[�GU��l�������	���Q
kGUQ���Bm[��g�`M֧qG���Q�b����<��G����r��䶎t�/��I�9�� �|h�b�o��M��鯄xJXĂ�h��}M*ە�q��!Nc�[�	��T�p�����&� ��f���D���ȐD)4)��c�/�EB`�C�Ҷ��9M.�%6�Ѧ8N�&�D���b���1e��<���N���TĿ(�tŬ��(��]6�."=���UO�⋔߆)T9�f	��~n�|Y�I���Ur�ݎ�5��1���)XƝQ"6H@}ɤ�QV� �rG��U��6��)���z����̑���)b X����o6�&�šĳ� �<LO�_��k"�I ��{,�(�p�����Ry���`N��k����%V����T��?h��f]���C��b�i���~�$@u�)Q]�>�X�� �/U�8�j� � p� �h�5�\l:��(4:�U:#HcR��6>�Q<��`-j+~]f2>a|��+E�>��)��7K_̾j�Z�_pw'pA�����*HH�9g�s��!��rJ���j���b�������a:ؚ�t��(������$����_�5w	?E�9Q��/b�/L�:bɤ��]����͂��q>�
Y�� ؓ�6��{h�)/H(�\��4���}�)I�r�E��jNCa1���%U����� a�J2_<ɍ6�����\*����AT� Ҵ(�u�[ l|HS������k�°����樬�w%����]"t3zCԛB���k�����]C��k�D��{�h�%MOH��}�Z�D��K}�p<:�?�W/v��@Z���ݥ�ʯȰ�ډ�k��b!u:'��S��������no(����K�듧P=����K��o���{�/[�iF< � MĦl6�+�>T{M��G8 St���TX�0C۟p�T�_w�+#���ӂf�jyrH�퍓G^�%�2��* <J�
���mW�\U+���[���P̺���0� ��F���T�k�x�X���9&B	��ݘB��Q/����u�z�S�h�Z��o ^����c��1����C0�ic�J��1w�oQ~��@R��A�A���!����P��D@r膡��A�$���PZb�������u�Ŏ���\k]k��j+��Q��MS�ɝ�o/`��h�2�T����R��D���ԏ�^�>y$gݴqk54ɹ��hY�XxϺ<,-�c�g��$���%�Η2��c��i�'��$h�D��y.@k[��GqM�X� �C��6�-�p�x��$��Ӄ׿��i��_�L2Q%LѴB�".uG�)�5T?�x�U�,�m��U�M���on�zP˕��342���hNWV�'}.z��$y6yN��y�EȐX]�(��4��W�,�����|���XW�R
�루# ��Kc�["ղ���,Ǹ?�����7�܌�i/�ˇhE�?��l�"��??�]f�'�/�ydTNX���/͢�o;��f�m�{¬���W��ӧw��mfk|�फ़�U��J[�H? ;� u��'p	��Յ~V��>Et��>Wx�ϙ�^��{Q�gu_a����VBTع*QX�¸�(���,եSApSp�o|5�Qè��8��3]E=P���!����!x�ft�l�{�r�_)��:9[N\\�+Fٛ����Y$���u'�3a�ank�(7�;=bd��@�������8&�ޓ/ #�=�{0^#���;Ŋ�g1���WMnzx,�����5�׉Ȩ%��8��v�C��7�]9���.�����	�לs��۔8�gރL<�k٨�5���s�H�"D��s~�<�S�fj��#4�&��b��ulfex-\��E#NSʿ�N�A%�g.��iu}��R��wW{Uy�=�"tC�]Ae�A�rwD�}2���y P}ҡ�>d�U?���̩
������uK+XO�/��X���d\&GԿ�bOrg:��Xv���Y�B�}�`��Ec�m�X�њN��s��v����3Z�,pʍon���[xz�H�kw���rQ�� �_����#�N�9��wԢBA<�o��vn>̀d��B��[z�W���թ
�$`��yL��+I-aѭ�[��xO>��U�85p����J;/�_�&��^��A��F���8MQ�_��Sך�� ��5�O�B �S���&~�ex�D��`8yp|�^k� cF��/�=$���sF��IqJ�ju����~��W	'0B��H�vLee��6�|k[��v�;R�G�"����#��sl��TIo��D@����͛��S2��
h���bt��j��F]0��>�C��T�Tqw���Yn���G�dD���:}� <q���~ͦ��/�Ea��c�޺%k��x3޹��%���R��f(`�Am�i�b��r4��

�)�VA �+�Z�D��u+1T�yp��l�nc��1���# �=R�N!����0��a��ޠ��(9�o��6��+w�=�Ox��K��ʑReG4%i^��ǧ��Py(���L[ ��/n��O�wE��O7�H!.��/]��h�t��?��#&����?��������R��,��8� -iF�_�Wo6�q�\��z���y����g����x )�X�}�?�L��?�� rӔm�2��bs�xW��	eA�f�C�&^���F�L� �J��8Yȡ��4�A������$G�hzDz�]����!��o@	N��ڳ�r����O�EƎZ��~�N�i$�xs��`ĕ�&�&��a�B����a	�ymbK[�����XEѣ�s;64V�bQ�y���/�gX��E_+�:O%��  U�l�P��1?�	���Hս���� }�2݉]���iu���ʯɾ���:���cv�}><��[U%�A�����p�ݸ��A�i��0Z�f�\̝���r*'�{?æ��%��F
bT��*�B��������A�M'�bd؈������A�+x��!=.Cܪ0�%�wH�E����׵͙�����+����������LIL�i�=;I@@p�����D
pY0�X�^)0Ƹ!�Q��]������+�92RY<�I\>�jzs01C*��z�㩰§�9y�M�[�r^@}�Gӎ��}.ʲy��ut�%`b�kx �F��L�'�a�g� x�Փ�ҷL_��R 5���tZV���}K?��՝\K��ܗ��p��:�|���X�&{|D��l
 �[�T�Wm5��&f�Q�r'��/^��_��)u�դ�)|�Y=u���S�~ �Q�"��;����?��%x���{��ɭpS��������
��Y��d�>5 !����"ʳ�w�͚mL�H�$��w(Mb�����Q��?/N^>=��W--�ʹu�ύp�zs7Tڂ~Jf������l��"�Om��䇩���r\�9��i�
�l��W��W�G�[Ed�X;g�=�W�?�%��U�������NR���wq:b��-͒,�m��$ghq���6c�@�Oܖ�>�{<����i��W�f��RӜ�������i����ӪZǻ�����Z�J�(\���������$V���	fz�2����rわM'��x���0[jFht�|zΖ݆��@�zD���AoG���2ZO��-M5�_�u��=_f5Ǘ�y B��m�*PK�,�+��K�.���ΰy���Fj������ػ����3e�|e����f�f/�_�)��!d� �l��Wg��I�س����?5Ll`�P��[W�##�6�`�K.RI��L��C<%��\���������K�m``r;4m.��Xk�Hp�J��1�-@o�ɝ3�TR�4�����z;�I2:�W��^'"�oT�$��.pݸSN�"߇Duao��Q���4�U#Ӗ� 9�{��Mߞ�d��ֶU����t�kY]�Zċ5g�����C��t�ժ�ȣZlfw؋6EB���͛Ep��t�+�x@����kzǮ�+S	��xf)łO558G4�;�2Y�S?� ��V֒�)���Tg��3�.�;�F�A������K�&�G�MAy�����̎���i�``��\Qz��lAhя,�A�,���V�`y��P��m�����������u�\� Y��U6f*��0l-4��:��V&ݳ8s:&wAmR�ȾSsQ�S��\�T;M����Y�2��';m�R�L�;U;I���	"TZ]R[�c�{��~��4�̈́
_Y�i^�`aF>�i�m�Vp
���Y�]+�
�W�`n�\�čG�X[C����h�Z��|%ߛi�	M�=�#���_���}��.T׹����C��D&����r����]�Ns��p�?oS4�������Gn��ˋÝ=�)$(�	�8j���i� �n��,ؖO�T��T��V@,�YB[�\����S��f��5���.�պ�&R̃)���
*c����D�%� S�.ꉑ,,�Xx�o��S��K�~�:��v�ok�����讦�ݸ���9?l\��b�x[-�����laIΩ�� ��~PW�2������A�u���}��C��;�$����67g�ܯb��Ř�7��V�"�9K��>m�9�-i*��%��Ą�2�̅l���/9j/F�~g�̦̽s1��-�w���]!����<�"�������U�B�Ic����-��_�{��Eǘ���j�PgE3���g����]�O�ﱜ�b�Y��w�>��`��k&�,Ȃ6�"���{�e��L�{r��e��Au>jM�pT�wҭ�2���p��A����S���^��O�n	��cb�q�ghW~�J�-��E�ך}�/s�o�!MH7��͂���Q�����������#�,�~�1�����b��^�zl�e"Gɨ�HۚS�s|����5G~mhk��H+b��F�x�
���d1��:�e$^Q�m��Y�C[Pz��s׮�]ю5��(�]����a�L�4_�<����$?R-�dxI�NX��� ��3�Q��Ʀ��&%�v]Z�恽�����yen�+��h]1�q %ن	K�ټG���>wn�P��*�{�S��L�gu��8o-�p�|'��k̒c�T&����p&4Y�F8�\��3�C���1�A]_�T;������d϶)��]����:�{/���b�U����E��\L1��:�Zq�~���P�26f��܉��)���5De|�U`��G����s�Ck�[bEC$�,񂸹`�oӚd��K���jg'ޟgT����C0�qr[���M(�(�<r�Za��R@J��F}9��^��l�#������
��m����'�{�_d	/e;�ǂy���$���V��߭��G@^R<�8��j�|z�	D�̸�/��Kl���}��D'�p���/"2}&9��Ov�q7�
|&_ 8=��|mlW}D�#�Ő���eei<�3�u%˗��1/�?�a���K��̟��'&����T���gF�Ι�m�� űT8�� "�H�i���t�o'L�V'/��X��Z:,��#d�iV.��K��@�Y:xd*bb�H3S����c�M�F@@���O ��Gd��|��)}��r����V�y��?7t�(U�z F9����,f���������{�󥆶�}���̬ ��9�#LE�󣲖քX7�ma��+%�{�'�}u��^��iV^rv��������M��4��8��7��W�>{Y�C-)���˴�$Y�4��Ĵ%PM���in=8��֚��*�YTPYqE¡����ե�#V�[|�I��?c���7��|1��d��x�S��wa��+84��LD�ƶ�o�e��T;v��I�����.����u�+�~�(W��J�|�z�.��&�9k�m[X=�	�P�5�䅅MTk�����O�|��巈�^��}����t޷Tx�WE1����ʠ����g'/�e�F�b"�1�J��c�e����I�\���n�e	M�N�IװY�J0������2vŰ*P��A�SN:�l�d�!�VS��<6��y3*19�%O��$��e�����Ӌ�&�v�hrIʓ�R�룅��v��ڏV}�X	1s�I��%�Y�/L;$O�# �:0�l))��DJ-���@�mo��ɸie�����qS�$殽������l=~(>_�X��Ēp�+x#���ba��Y&Y`e�T�������4�2��}*P��A&�#�V��R�1�E�����0H�l��M��O�ރ�P/���{�l�X!�"��d	�b;0�s�q�g��U�J��R��������t=��2��KUd;'�Ɣ��g�*�3�܀6ʛ�D�S���gF�vq�x�,ި�g.e�on������Y��c�"*�r��Y2b�<Uԛ�|O(f38&d	�3�OG�S��ؽ�7�b
tNB�)>g��y& �ă�Pt�RLq��br�L5�|���uv�M���6��t�N۞�SK�*�;��s����|�����x��}�U'��>����vq�n�aʃ�ll�=�t�0��L���7(V-$vo���8X��-&���37��Os=W�!�N/=X�-hQ�-�aͳ���HwIv33�������0��Z������d��OM�n�bl�I��٘��:�S�Vo�jnU�=
�FIt\�u�l�F)�
��qE-d\dS:��Ϙ��pK�2�I!�%A�:c��]�Uz&2��HONk��h��,���,�7�d�/?�Ӕ����`�xE�_Wg�a�pNkJ���cq����?�x���rV���;�����㤎�'��3Ȣ���Gl7�O�����I���G�|{�>�9R�S|$��`H�s�ӟ�Ο>�Y��V �Ē�fY��y�4���)�����@�0�����C�q|��K���&e������=~nt�����e���q�����g0�P��-�D���Si���ݞ��y�Bm�-�g�/9[�������0&�+��-u��ğ�8�16`��~`�b�_�^
>-0^?ػ&J�7m���ȿ�j�0�/[��xȤիG��]6�v��;!GG&�ѩ�	�������@����au�������	P���sk���p�tTEM�Gڗ]2�ťj�`D��c'��_:�l��z�`V����#s��^�c^(��	�a�T6�6;ٚ���߾���3�T=}Z���V�����0}������/�~�U,��R@�B�I����ߤ��f�E�a��7>l�����F�l?� 5VؤxM�C��mU��K�­өų��%Lۉ�)(� ��0+����U�8�e�У�Z#۲�|�j��}&�0f�����&αSQԤF09���܇_��tߏ���mݍ/�
�(r��
�x_p�|����.�.9۩}ߔ\�w��C�8��}���V��\�Dh�0�N�����x9.톲�;�c>�e�od�C,���S��\�S��,d���S��;0x|���qA�x!!��;	�n��a89j1���(����W�U�I��l��%����}z�A�^�Rs�����n9gxZ ދܙ��wźP��߻8��&�<�oU�����p��7u�Y�h|��O�4˅�`�k{0�힌;�:ě��!��7�kD�ew|q��f�c>����
>�c1vW*����J|�����o�ѿ���3��j�WN�˷�P}�ov4���Ñ��9���$�@�be�gZԈ40��!�ǵ\����)h0fyI{�����X!3��U��:��׷��ђ3�r�5P�-����H��qq�`D�2�3���`�����ڦ#�,+K���S^�Cj�0(�j%C��1�|)���f���Y|�v����?kn6��>F�rFVHT�<P�� �&j]�M�7�˻��,f��g�m��<R��jJb_I�I��&S7�?)��6�6��e3����?!���!0����Nrrqɢ��Vޅd(��7E���+	�~�Y�D��2�oc�^F��O��A�[ل�Db���g�:������aQē�؊��d ֋M�=��:�K�e�ꇼUGҒ���Jً�y�0F���o,��4��B���ȿm>�U���H�땐H%0I�F7��z����Y�"���{�x}��x��_�E$���r��F���$��K���{L����7�]��`�Sn�������Q/�� L`D���i�~Pc��V��2%b���q@��Ʒh^�h�	�FX�X�
��Nw�[{�k<�a�� ��ڕ<߸��8��-t����=���������#˥2��Bo*�<����9�=@#�2��A��,�?�s6�\RҢ|�*�K���0B��2��d����x��5�����M��'��f��Lݠ4�*�+!��.mL�0�25�:*>:t����T`Ƚ��i�ҿ�:��9Ս��C�Ya���q�2H�`��k��Ղ�7y��=#�#m^�!��2����V �ЈI� �� �_{K�%򅣈h����R�F���$qD�/��w��s�g���hz�(S��bp����Wo�)���Q��p�_r�f�OTߑW+���ń�4$��&Hw���\+8F�t&�N���o��%>�W-���!|.�+M���7��hnȈ���|�CD�l��e3:�\4[����Ļ�kES�b(S��"�]�i�?�PErd��qڗtg��t�Ti!��FG1[�����0-M��>d�m�T?�v�ೃ�SJ�]�ڧv&����
ȋ�+�l墢����yk��2�D����$��{����Z�}^�g7��Q�a7��9��!�6�_�XS ಾr��=��<1��J�)#�\������-�(	����j��ո�����:�-+�R�QN���:3��Q���v�
n��/��(S|?Y�~ Å]ALRq���:�ra���AT}���1GLM�FwI���	iR��l5�ʓ�}$;�&�
r���W{�5����}3s��r5��g��3ޓ;��<smrr�ӉB\S��H���qeH<7�ϣ'9��/��y�*�h���,?��#½�-��޶����߁��#&���O��;�g"���?��M	��O$��@��&Kſ��$���W�g8n�r3��wdO�VD��+�H%����^?)��0GZh����6Vw"��m5wg�{�p
�_1+���~������ ��|��6��_��K��2�ET_���^��誫i��K�	���x7O�)�m��P }
$�����;+k��h?/�����ݚ��`A��Ĉ���"di\�������'R���%ֶ0�z��C�ܟ�/ΐ���MQtxR�R�~a���%٧L���8B�����9��;	7xu���>�������}�R��#@�V23�Xw�e�+�ͅ&s�~?C�ճq� r�QR�'�����۽�:K��앓���X�#3p|o_EzMm1��$)4K.^C&��z�2f˝����GƐ{)+z����u��L_#��#�����2��:�e�F>��>��fv(���vbT�g%w�qBB"�d�2;�=�v��N� �ۮ*�\�+x$L]`4�nu��x�A���+�T�3-L�u$=��(��֯�88�.�eU��8:�
g�J<��yݷ����;
gs��/�Z(�:�θp�1�%J��_1�7�l�%kf+�#��F�er�\Ɍ�z8��bC�g�8�������O:[�@�
�v-��k��/J&-�-Ǔ�_��T����9bs�E$�M������V��%&nW�:6�H5 �U��/du�<i�~8*@$�PJ�wS��~��35����R��8�%PA]E��3'�Ax��Y�xW�蒾	V��*Ȼ�0�m]�r�ܾ���[2�E�heN�9O�,�@�G�<=�b{`���Xk��o���aM�C�M]�Xq�R�j%�����k�5-��5�s�%����EҶ�)�����:�hf�j����R�y��d�F���ɒ_�R�����O �	���vA�zZǽ8��lY+>�:����%�	�94UP̹§����di2���9��G�뗜���B}��nj�L� Z�/�>������d��,�d�3'��y������S���t8�5O
b���?���nG3}��8�H��A� R�dp74��K��ɾ���8W��۵Ք̣�\N��ݳ����/:m���%S1���L�R���\r���kKHS^�gy��{۪�����F����Q�qCy��w�����D�e2�^�Z��9Ef���r�MX/ve񘂫�;�����}	��_8��Wzvd�����+�Y��r�1Ε��U��]@zWф)5.�����7ϻ*�X,�*-��@�#��ߜ��7�Pt��ZbΉ�a�a�U��(�S��>x�w�̓���Czۘ&���R�s�~��p�H�(;�{��E���R���Yʑ�>�3Ʉ�?�}�"#|�o�WV�.�-��z�J���<0�ѯ�e���\p�����ݷJ��;����T	�gW�����Ύ�w�����[��!�s��l�F�։�ox\����+Y݇����M���������r��i��'c1�X���Z����Θ�R���O��p(I��E�Z� C�OC���Bl��
C����Q#6|�o|;9vs��{I�I5 � \uf-�~���koB� 6 �rc&��'��������2y���[���D7Z�)ŒԱ�?�8�?*LZtt]���C4��GL��?.>��M5O���+YY�"�����"��ӂ��d$ߢ��j:V4�%3^��uB.��J�� ����0�m�B��_r�,dn"_|��,@)�ap�ߞb>P���q�W�L��!+�95Xp �� z�=���!�$Zp��=�t��q�@˓�O�c�����.8w��q�:ԍzv�?:jޅR�XɕU/Q� x~u@�(���5|���b�d�\�F��)�7R$�3���A�������:���V���kܛf�U+�4ZC8�8���V
��Kts:}x��n�}������oo�_^�&x	~�S�ޡ"+��?ÿ��F�|>��8���i����F������hoK��by��qx&@y6�;��f�֌`K}����!�C._��7��0K, {�-�yG���bL܀?*77u��Y:�`|���(�[�,\���&"��c#q��&ee:DR��'%�֓��Ά啚��K�6 <��)K��i��-��&�Z�H�	BZj��GԫzG�'��X��^�^)�b`��C�e��`���u���	.×G���G��yF>��MT������H��>^�^F� ��zVeS�HA����L`��k��:	��&�kΕ��޾X�:L����b�/4X��E�8��G�d��+$��A�pE�zpm��)��&���*��W?���~��sc�p+l�!���N�w%��l$ᓼ���8�c�������9 ����\F��<�~h�}��c�g
Cy�u���V����/v���J2�ڰ~��iX0��-5�0������N�=\����\�e��h\@n�_�5`8P�����3�Fb+�N������+Pn��V�U��r�tX���6��v����aƥ�mM�?:�4C4��\�FV�w�ޛ����(��%Hh��}��H\7�'�F�s�$7LG�Y��vJ�W质���N��U������%O���3��ô\B�-"؅��`j�����o����������P��8T�+1W�����v���I�2���������{ =r�:w�.߸�y�1����Gy�A�+>�;��a
6�.��*�1_�X���C?;�Y�:u�*���6��]�zg��0��3ru�w2f`w2�hU](9�����d����E��A����Qp����I]���5�+�Nc��gMT�2Cƾ�e<I��b��v�&Ar�>�yXK3���*�3.=��٭��?/�� 9�ݬ�{d��x&�g�O:�Ϙ8s��Ң��_~��0�ح+d$(�>�E�<_�L�iH��@�bC�I\��q���h��J�_E����n3��(����f���W�:����s��Kv�vV�s'_��:���n���M���8;�XL0��`���[�������z�+�i�ϠG^g�/=C�B���u�����{3�h��0�D�MT}�K�eB��,��"n�(�g��z�7Y��gF�$�B¹6M\B/�vp����@���������SίO)䜍���D	C��������>��J=*��hY4yy���b�ָ�����
��ڹƵ�;�����e%�����~�;s�?K��H
��i��L;�ə-"_�q�͝�-���X�zYΪD<��w� G����$_���ѫ#�Ծ�k$M��-V����޿+��Yr	f�ݝtw���~�R1b�A���h^�]�GS�{F'����a��F��,�V������H�v��T;bl��pe:�W��˗��ǎ��ъw�˸f*�驰�L�� �ď�p�剣����O�d��Ԇ�J�����5�@��B�η��'uh�b�Y�=�ݕTl�0?&���|V��_�Q��}Q�l`�׹�[�Q���%Q�w�\�# �\��K�8�c�.�;!�q��"�X8��u߈,a�[������<�/N�֒C�1��]?�\r�$��5��]���Q�gx*n��/���r��oY@�v�;�!O�9����xAIb<ǽ�ǜa��\�j�&b���TN������Ʉ���e1��u����e=��Mٛ쐳hM1C�Jp���k
�剗WˢW3?�Oޞ>��,d'�/��Ӻ�{4�|q�5���R�����u���F/y�����Z�A�\t��%��X��ݰc��Ђ?��ӵg�o�'.}��m�/}�P�������rKq̤&������{9�/)�fyq-[�gse����@����-T�Bڟ�޿�`��a���K08I{�=߆|�ky-�P��z������M'e!֋���]b��^wl7��P�Y�or�ڧ����o��w�lT΃�$��ԯce!k�0ؤ��T���i�_��Н s���N���?�b!Fq�;�H�cʕ��Pl�������]���Uø�!���n&�%�܎/��g�N��&&�/��W�T@Tc��t�Ξa�;'��5X��`��@�x\��̆.lwſ��t���}�;��;�s~h;"��p-Y��Iin��l�/��w{�K�=��8lxPZu�{�W�'����B�*~�hx*VQa�o�D����n{�,�y��kʌ�qO<m6�^ig�v��C:����ԠS�|�/�~R���?����+X�M���ٺLX!pL#��{j�qOur��%�U�Y��
�'R}µ�
oS�N#�;���̃�yE�l}�e��LEN��X(���F�x�q��G�O�������=�e¢C�
�k5`p����wEjGN�D�b��W^�aF�T)J����ϔC*`�Q�gmV�Q��ϻ׫��S\�b��'˦u?_`��a����䔇�l)�=���<�����9�*��l-ծ���`�a�s^āYe����ɬ��	x?��["�E�C��"
	zpY�q�V��J���n[.���S1R�-�8yov 7�U��z/���4���"�с�U5J�e==?'w#�>�����]2|E��x�Q�/��3m�3L�t�cu���W�Þܮ��-��t��Er.=�w�k�aIg�s�]+�邀*�ΣB�l4.hv@~W,L${'5����'��f���x)ߵ��)�i�3C�}��qs-b~�19g'י�N�6��HK���M�pt��U��k�ĘQ/������V_���Iz����%|���B57��\���E�����<�yˍ��>�Ე��.C���_�3���o��r���|%2�P�8d�0��Ѹ����֙)>0x�}������#_��J�1v��%�T�8�W�\C#@�л��+�l��#��aYE[uR���`̥���|�.�qoG�G!�XQ���E�4���������#���#@�b~r�/����<F�Y�b��B&w�w���·@�E<�[W�٫V�����7��B�큾c�x���4���%P��9_��C�R���U'EE��q��#�T6
�H6n4��.�F2+�$�.�lT�O[gg⬼i.XU�1���LH�嘖�oX�9�D�>\Qò�A�?e���q������-╀:q��-�D���ᄞ�]j�t�� �G�9F��a*d��1�-�����J�8ղw�M��A҈���c:L�����b�/q����yl�;_ٺ���V騖X�aEz�:Yh
��ǈqLmN��2}�'���9�ǖa�v~{�wq��/�����|��j��R	�9�8?P��0�$,�	DxQ��ڒ�J7h����T)�srp�8vS1qz��W�d��%1ZYJ� l�U#�m��P�����(#Ŀ�o�y��b��(ڱϽ���~�]��<�`�*Y��^��S��"v�s��#��p�9\͖�Y��T} Qi�Z\�IFHg��$x5W��5�%0��ҫ�I����F��9Of>�'�R@�.��O��F.Lii��^*T����%��@�O�"4*�u��H�j/�%b�j�l\��D��������?���ݏ3�'��j���n��̬_���,.���
����d
�sC����A��"�/Ԓ-�]�ţn���E1�J�eFu���LĬ��l	�_(�����Ȳ�Q���6����Kh�v�*��r���a��n�T� �����[��Y�=^��U,���r���Ed�u��r�A�����i)$��h��=)e���	�?�k����$��ψ�Q�{ �޽h�FS�M܆�j.J��=T�_���[S#��3�(ŅV�B�����J�8X��������gr�mb�1��N��	h�Mn'-[;�ZSt{�n�V��1l��6�.�rhyB}��n�g8��K�[�7���&�W�ܸ ��c����c��m ����� �F�� F�L�N��ﴓ�8����2���ǰ��� ��O��Z�K��ͺ]�c�ն06tp�#KJ�49ə��wj�\
��0�)�/|[H~i��o�Ψr�,�ޝd�6��@g�DU�����lRM�?��
���H-��eM|��M���
��9����%M�ף:oE����=��/~6Ӱ�e9�f��V�o��b
gXh����J��%�F��iiD_g4��.�SL٘��QHtº��֬ߛ^Xb)3ƛ�<��x��v����~���~�����~OZ~�9�R�k�QpW�?��nW|��v:��q��o��΅uk����b�kQPh�X?�Y�A��`��*ܛ���_���*#7F��ڀ�S/{��L�6��r�<|NOZ ��)��2��8~�P�r��	�� ���KlJ4�j�����?�S��K�yB-��d��MR�C+lf�y��ǭ��6ol`����$�� Y禶�c�̬��Mcn�榪���`��ʑ���V����k�r�T�",:�Z���	@��ܓk�D��0���d�7�%����ʴ�����kRdVRw�y \�F-]�թ>%�^�B�I�s�/)�l�}����<�Ԋѣ�k��jx��s����Z�.��k����@�C�x��cŁV�iE���G�����P!lse���3�|�͓ z����(Y)��is�ޔ�5r�mC�{����U�+=LRս�P
� ��@�N��V8�Ĉ���a~P����P{��0�#�%�ib��Ś���Lm���L!Uq��O`�8"Nt�S Ԡ�,F��q��q��%5/�K���N�ӯ:������?%�i9���?F*.>

^���f���c�$Q3)(P�E��||��Ŗ�I�(�"�0��1�+`<O�|f,Ob�����|�(�h5Bo1`���l^�\=�����]���/f����$�(ܾ+)�0��@Ɗwu�ճ�����russ���tBA�T�" V�Ed�c٢,+4/�1pmP�/*<�h�л�c?�'��wc>jc7��[����A�,q ���@�\co���#A�,����?�,��eEr��L��<O狉[�9_�^\+���&*#�>����5f&I+�eX���`w�ꪼ��gfP .a���g�f�.��B�.I�D��i�N�1G��sW����J�Ƀ��د�*h��Q��2��0�좡g�;N�`�Fj��x�p�~�A@B\��㾻�RVt�b��O����4��5��q��H��c���m�G@�e�#`^7����d!�[g��r/8���!�AU|8qO� ��I��ØRm�>s������iG�2������WłB�u+����b��Zi�I�T�N�yQ���O�>�sC�����F�`�7$u��&��1�������,��|��(�<>��a�ۨ���ӧ���>:��G��?H��ɗ^/������I0��~��׋��s�nc
F}� �+�θs�͕#a��yA��^qIS�j�}>a�-1I��?�R�(:�a�3!���Z(�Ti��Yχ�p��$�$~
����Ѻ��eM��f5��D{���3yc9xIަYUL��~S��PkU��Ɲ}���X�п�М�$2��Ҹ�;6ͩ��_}dƋ%��/ǿ\53���k��x��x;/5R%��wg�J>#�mُ|k3S�c����>΢E�d»i�<4O�Dۓ�1�ڥ��h�I��w��I��5'_be�>���['�o73-�����yg�����s�� �63,?�^���~* �vG��"A�(���\�g᪝c�[��L}�Ħ����d]�O3~���u����k�awt��3{W�qk��6�g���QZ���9f�8�u�t�߱�U���6�%�_
�ٜ���Ϊ�yV@�C<}π�Quo���dj�L5��z8���:���W�8w���+?���D�!���u�]4�N��s�$>�۰v����s��x�D1ӵj������1�l�����3fF�`4�E��ܒ;���?��N�dن�Re�VcoK- }�'�Nŝ`��2U��l&�G���H�]��!�Œ�������:��hT���ED�4�/����m̛If�'S��
y�ͅ��OkMċ
�0ɩ7>��2}�/�N�A�E4���f�0�ĥ�e�-O>�����7�?��J��F(E���x�~eh)�pd�[<s(��\D`=���ُ �lg��EF�/�@^&��`q�n�Kެ��+~~�����B��k�����W��,��!X�Cp� A���Np	>Hpw��w�$��:�wn���p�=���k���zuWq�I՜[��h�#\�y����+��_͙.2�;�� �4CuNy�\f������GR`�G�C�̚لf�v��kR9<3�	�[�e��/��)�w�.��y��	
A���EZE���IBݶ��xq�ja��2��@��f[����Py츁���?�,�}p�x�r�Q:+�dQ�~�)��;\�Zǥ���Vxg�%.i:^�&�S�
��sϥ�rћ���)��������)HI0Q�{[�wrۘ��WB��{�Yֳ��N�)&���x���笇�eO*�.<�v�i�iZ����/��9e	L	D��fݭ��[�ߨ6�|�J�)��?\_=��[��~�l���R5p���~F��˄4tg���5w���w]��~���$C���9,_��X�����{#G�~U��WM9��tsɛ�b"�\\���1�\�H����Q u��-ܣ�~f��-��c�3�%�����`�M���������7���V��T�K˞�:�A�^	�G1$q60M���|�1�D?��w#�IW�I2n���.�C��WW	��������Q����=�c���:Y�
��RI�L�ÿ�զ��D��FH?�S�%��TW�������;e��2�}5�i����s��$	i����}נ�֛D�;���Я+_�1"���-]Qkg�`0B���+��隊(�N����)eyZ>j#������bx�"�;�.��_�w8�x	P�	\+�w�/�M;}�C�U KD)�û���R~���C���娏#�-�⠚}}�եU�"F��!N����@�|��^�����Xv��ZH��~э/WF�`BE�X�G�}nD�Wz|"�PJ��\������cb8YE������������0"5=�D[;��y{�(�{�V���hΤ]���ZX��aڳ��/�V��+9T�#�T�R��E��XI|<��z�}��z9��=�o�l���ݐD�k����`����OI}-;uM���A�	�L��Y�ȔX��EjZ����/*"+{\�-}�׸���	m���|�u�%N/e�1L�;���,��Q���*�d����9�W9����F���c�x��3�߰ pr��hk,~�m�@1q�Vy��	�' ���˿���Kk��p�]U_���Ŀ7�"���CF?��rf�rf9	�D��Y���c��8�V:%e���I�H�c2�S�y)R��F�{���K�����u�e"��~ZJ�6�;��G|��t�Χu�4�������	�И�D�x�H�%_t�<�˜�&�������i�W�G����m7�w��q��������� s��s�����*�/+?7Tf��Y���R�}l
���]Z��+�&W�3g�6��b�T�`2έ�dr)�q^?H�KM�ݶz�P��)HP��3I^�2}$X+����	��F��������]��=��f�d|�b�LtK̢��q�8�)��y�^�(Ť��G$����O���L'UC1A�����cV��1by�w�����s�
���`��h��@��O�'O`R����t�܌K��B�H�j3W�Ǆ3�p|jQ� -���П�X��R����@m�V���板��wA�M�W��v5���_d�n��Ѽ�2��� �1K܊*^�pӅ�̷W T����)+~�v]���}a}�10�i(Q[-rJMᠯI�S�z�}h�L�ỉ���d}�β�&V�������h�F��?�e��j�b�PA0��Ѷ.�V����r�-�4bJ�@s ��y�����|Kx���6e:A�vXU�=a����%+��VTL���W߯ �������``h3ee�{�v�"dIPR����	?d刘���0�1��#��6�� �
k��h�ɯ�i�˘F�7VK���E�q#Rtz�t��j��kc�%�T�j�6.�������JZT �X������~P�{�xuc}��P�+3$j��i2H�z�}$�Th˛�Ю.*��7�E���%tk�	��Tg�-��>��*~�!��	��Ѽ�)��l}s=~Њ4!z�QWU!W��
��U���k����@�*�7�.�Ōb������T�����њ|Z�ݝ5=��"Cx�Ԇ�\�@&�8��cy���n��  ��VX�k�����m��ͣsV��*�/)`	�ΎW�����.M~�K��-��'����L����l�����z�%Ϯn6KWH	���Y�Xl��^��g�v>�k��[ȓ���]��8�eCDS������~�hY��,�����{"2B�Q����Q���9:&Ǎ�ӛ�¦Ļ,X��+�ɹ%p�ͼ�W|�Gq����e�w��|��O�C��V`T�an�ݑБ���C���_HF��n��oN=��z����T7��_�M��Ы�K����+i9����Ġ/�
	)���;���c��7�C��Γ�����#eSD5y�T2;Lv\�|9�4"��ȁ�/���uG�G���>�iQ����}����&<]ᶔ�bV�y��&7g E�)�-}_�;�v��p�{��*���W���h�E���T�����I�%����16�,�g��$�$-���c��BC^�(ܻ$a���"�h��=-��.�pJ~��u:g'��L�,{oǬ��)JR"t�v8_�	��	�%��Q�u'G�԰���C��#�|��7ej%����7��� �":~&���9)1�s"��Ǜ�r��8��S�_^�ӄ���
��j����B{���C�0+��'Ww�;{�4ٌ($ϯ����a����U?�&܆F�K�R2qL��HV�/��0W%=1�2�:���TQ�����M�{[���
�[�Y�({7%��[it��cf�oT'�D�/�0��\L�{wR9��F'>����&����:�׼�̰��?R�Y���P����~�x��#I��{�em��(�b?��7^Fs=�b�Λ~�J���׳�ªO��b�[{*�J���wbO�WifU��@a"������[�yG�7"<�[i����A������1�B��3�SE���ؤ:�͑Y%$�<�s:�k��j��@��
@j��t�,ttն�jn�~8",	�Q���q�>�ʓ��O��^T&����i���b��ީ`�s���;�n��J���� A�H=�p{�\=u�7T����ɝ����4A��zW�9�v@SJ�͠l]�cy�s�n�a��vN��W;3��^!I:i	��Q�V�$�զ���v�E=����S�k��Xn�l?z���	��Y��eD&��.����g��W�Ej��f0Kk=�?�;~��7��3��k��#�͗�Cߠ�)�
;/w�Py�呈2�3�A��D}�Q�G��C��~cR���S��љ�\�&���
�F����bq�#y��k��H����ܹ��$����?	b�;T𱅝���D�CZ)ʖ'C���/A�S�����������J��Jfpaּ��.�\�m����P������ýM��g�䉯6_T��E��y� ���<�_>��$Gu��#T=��ʩ ?�Qήu�ǲ2ƣ�2�p�m�ō�n^V�lŔc�Xk�;} Q	��aDnꁝhd�><,D��g��	�x�����%?*��XV'&��Q 'wP-�p�C�ol4p�����-i0�+��+ fR"�T�1�p�,(��ǣ�o?��K7�7Z�f6���k���l���qv!?.9���9B{���/�
���W[�!�pn��y�o
F&��[,P��9�=*�7�+漬�H�!tFv[�q�Mll��v �>�AZ���,?����W~�_������eClh�����-��@����	�M#ʇ;�L[�������p4Lj�/[o)�%a�u�@\Rt��Q��wЌ�t�o�<
Gà��e$��M&S�}HQ[Ng]��k�v^�7� m7�O8۽�8ڊ�d�j�R���)<�<��a�:�{���h��Rl����ąj/&Gi[�7I��n"�JtsH����L������IM���HH��KlL�_h����1�$29�M��������;w	��M�ť���	��!�F!�Kݏ!�a3�����d�6kr��_���WHE��#�L6���6���k�a֋��т���1mQ,���e}��d��9eio3��������R��!�1kh7��ƏT'g�e�96�6�;�܏�]ŨBy���
d�l��I'�ჺ{��f�-���'���U�j.U]�÷�ΘAg'<��M(�4鹛�4�zo�߾Uo�)��Sz>��!7��gZb-L�ՠ�/��Ŋ��Ļ�PY�R�}.�PQ��V��'�k� ���ı�ؾrE�j-���1<R�Q�UK]2�1Ȟ�I��m^�8��W1���4~��'7�(h2�&�'h3��Zq>>
9�~f�u����tC��������ѣ����������J��l�w�%���W�T	�_��(~<~3�DB8"",B�]\����r�ƪ�j�7��OiN�	���X8~�&����Ф������U�����8�[/<�%Py��Px�2z���$a-�������z}����r���')�Z�+g~u:~jؓ�϶#�c�OM*?�ȩ�e��Y�5]Fh�S��%m$�o:%���i�C!��sݞ�;���6xO�2�c5g\H��k�ΰ�r���v����d���ϓ?�j�ڭ�я�4�����ߩl�?��z{�\��R0������sE'�)�Dit=�=��w<��v������~�%��w�k�Nv�]�po��{�����(R��P�)�c��|�`�K��%_m8�Cj���s�4���Vסk�*b��v&�r���N����"����^��5�갰E"z���$����|n�
#����]�?C�ڠ0|����+��*�j9��A-������`R�t'�U
'�r��L���%���W��wl���W���W@���p�L��׵�`_���I�z����k�3PN�W��/���9�BR^%�qw;��{�����M��� �Z"~�{E��?��j~��Wo�=���\;-��E������R^�����R��n�>��P��
<ؾ�Ag�n2 A_�h���Y�ս��ߺk��[��C��8O����x ��=_�l��OX��姨���˲c
�������!Ae���� �V}��<P���|Yo�]��+f^-���4u�>���!$�Rԓ:Y�y~ZH���o��*<lP�/������/Ԓ����Zh9ss=����dG~U+�����4 ����}Q��>N-&�t�3<ܩ�>�&� @jҧ�AK��θ�6���|e���ܟ��'K��2��E�F�#M��c�!Q��5�L[�+����I�$b�|�,�9�^P5˳�)�x��NW�aJ��&��ٌ�p��yhC���\� �+�+��γ���ي<�7��Y۴�c��L��iP�0�(m��I���ˍ�R	���c9�F?��4,uX}I�A>w]Nx�4�,��7"��� �����[�H����]X�y�����w]�]}�V��$�aN}���Yy�)���9r�Ǿ���Η�޶�(`�xAٸ�����M�������\a�u���.G�U�����rɪ���G��8�����r��`��R8�����~���X��y��#�چ�]�;M,�Dҧ�}�]x�X�[���J&T~�c#�6�����N����}���x�� ~�����/@���è5��Ɨכ�f�Z��r<�<Og�d��ϸ4
3?lW�B�~ux��d��E"g��Cl���c䎻HSN˲q/��h>ki��as�,W$%h�*~x8��м�Cpf���$ɪ`	(d�|���ED��ڿeUQ���0��{�نՇ�.��M>љ���H��3%r�_��:�>�!���O�����9	����yj_�2��/y�{�
��X��Y9�R:'bI�XG\��Otɬ5f�G-�k?!���+b�T��H]���S��z8��Ϝe�b���&+Eg;��?唲q�c�|���Q���W�O���c�9���l/<����ݗ�UdY�23��D���
 CP��1svFP�	�|��K�\��>l��\)�/��r�e�lt�#����:ص��#q�`�s��i5�ְ	���`����7ORE;anT�l?:E#	�%aR�59l%#>(�⹂�L*�Ǉ�z��^����A]A�F�8)v��VL��}�1W<*2^���V��m��
�1�wMʼs��?+�610^nkB䞻�cY��9���y�ʩU�hd�Ff��a	8��w�_��ު�`����ܡ�U[s��|̰�LU'�"��P��P-
XP��x�Rv� ��;�Φ���\������4 v�':aB[�
�,���B�a)E�%Q�;��t-ck�F���_1;�{���xW_F�L�lw*X���c%H�cv�t����+K�Yw���v�P���ގ�-T8����j�?N�Yfz�� N�=��I���9(��]�:5J���0�|xVz$�$lW&j�;Z��;|h�]���@x�N4��e)��(%�{�I!-Ӛ�82権�����|��E
x����Y.$��U	5J��\�rq�b�g�k��ODJ�f�l /�-��u�9��F =�x�yo�@6{��o{�(l�V�ǅ��oj�;�����O+��.�7���_1�GI:�����#?�϶��h^��m�qZ�@�'n�)e!�� ����A# CMU�8/^xd�R�c�{�"[�@�S��@µל�O��O>����E�ٸ�F�8�.-���a��5 �NQkfP��͏첅��-T��.��\ �B�XTI�>����ʼ����w3Ԙ4�DHZ�M�"ҋ��Y��f�jq&�a��+ �1@�q��H���������G3�Vto:��� �l�j�WI.'�q�ZԠe�Ǉ�j{
,�1W�E��,򉨷��fl�{��]=��I��6r�(���#�+���}ZU��é�i��^��UTfv�G�˼��Kn��h���ܻ�݅�l�r�,=Z�9���(:wm�b�o��/����� w�`�=�$��Ql"U!U<P�*
m�r���f��%����K���F�zK[�9�f�E���<x���R���~K%�do�I�>r�tҭ�%��+	�_3����ʗ!�t��E.�fc��*��'&hY�_~;�M�&*o���[oY����������Q�Yl������
��Me��1�[��='������9�W6�4���	�Mxߠ뒪��$�C"�����T�W���³&1�q� 
�L�/�w����g/��_�Z�ZR���;�B�߾u���H�u�g���{���.��&��fbO�1��G5�AO��-u�,%��j�f*Hf�-1b����0\e����S�H:�
�����S��p��p��J�Z�EZ�0���ǱfIZ��t��Gٛ;;�R;��2e/�mMd�J�2i"�W|����2�!}}0:�*�K�AIo�;��ۉ�����+�q^J�N*�r*�!S$o��i'CN����y���;9��!�=��P$��U��h�Va����YU��%u�I�𴙛%�4�(n���<�|02��H�A����k&ؑ���c�����ȟ��򨻫j�Z�Ϯj����W&�"�ͥ�\��4B���߸h�?�%-��)^؟I�L66��$��B���|����#qFؤ�۾�}w�Qm*���Wf�?,P9[�	�Q�&� 'Ы�ck,5��0�C�Xڐ\�-I��K��:\\GG�B8$�\w'Z/兜�<ht{Zc��b2䏐�N3��Wn�\q;��H1��ƥ,G '��V���f�����2��賖^��Nq��?���Y��!.X��֫�G̘ 3��H��_$��Ǭ��XMQ͑Ĉ�h1rY�&��:�Zǋ����B�Gv���%�M�D������T�k �1]�EX�#Y��a�pk�i_(sy���RUM9���nVH��°&C��2&ҮÓ��D��y{Ĩ\Ա���S~��l��I��JA/FƑ��E���`�^����[9��s�NAnZ���_�������\��1�ʇ\�M0�@���,Gl�'�?+���F��{wk�nT$�/�-�4�:?�*v`9��l�8.������8�K��y	�Y��v���*�]�~�d���r	V��}U�ċ;��S G�0�cы蟅��b�	�{6�$-a8�����^Y���<�c�
�/77U��͙t��2�0|�P��j-�R�j���O�y��j�!�>��"�̼�wl���s3������##y�77w�l�3�A�,���P�|a��?����X��2���ĉ�K�99n/�����
f��Ɂ��,W�7�M���x�\�7�R��Չμ܆{�Z�~p������t�3�@��	�҉o��C<p�va��P?�
`��d�Zc��j�4�%FS�]��`nNk@R�C��g!���B��?h�+�'+�~@�w��H>y�ܰ<BQ�k�&@�����P~iհ�������YM���:�J���V�h����)8��\K�jLx�(2�%vdQ8�n���ҹ����t�ȅi��?ח�b�����N��݊$�3��PF.�8"Ͽ�fn�!'��5�B�E�KH�9�a}��}Fz~xm7!��]�v	=yx۱�r��6�T�l�4�Q:ve�Ck)Ni���))30V�����~�ѻ�<��o�
Pi���zpc,�px�渣�O�",�GB����iD�]M�c;K�a�K5�[ߠ�����҂�
8I����*�y%�^�%ۡZ[�r�����܀.Vh�!�QKæ����$����I=fH��s7b�'�=���?S<t��=Ы�9$�C����5�sv�ΐ���ꇽѿ�JU�A����H"��I���K"{��>�}l&�̆K������HRFe�7�o-��3��rc�f���Ôf"A_m1�s\iW^�®��m�~�Ua6vB�(�VNf �'�WB�V�����m��i������f5� ś���A6�Yz��ɏ�g�����j���-��r�Җt��]Né1�8�!t��XU��|�����~� �x@�Ls���(�ո����T�������y�S�b≒3�L��C�D���*�挂�w`����]*��榶h�R5��'&�zK~P��A&�����/���}~����}5|����c+��%8C �j���j�|i�=?��8�r�,�ِ3�9]�ս� �O@6��2J���kΥS	"��LRP%��!k�J��(Lz38;�L�Z/�jF�SO����!�y�[	��,#Y�݄�k�7Rw���p���[g�n�^lv�E-E� :�VD:�+ ���s�fBD��i��z�y�ܑ҅�c�;��"�$+m���_,@���Ew�&��Q�in@�ߐ��"��9��˪nfb��R��^�n�BS�ѓ�v\0���rj3��w)_��b���3$�YV�jD*:�B'��wE�_fd���:U�ڍJҿ��[�b��_"63�N˯�4~�<Ni�����d�LP]-��ZbC��Q؟2����4��u�PX+7��97eٮ
[��%j����}��kO�t?L�2�$�Eϵ��z1�~��t����̦��s��Y�D0�e�)�m���)���g��
�j�C�}�^�2Fz��E��g��ѿ��a�G_w�Y"0�%�ŕ0>1I!Lx�Elw��� S`(�EA/Xo��X%�KUqg��pGE��/�F��wE�==�.��W��2����it�51@�[�׵>��X����l��H���X]h�	����[��y�Բ�W9:�[�AeY��w�ٛ��|�y��{�� e�Om?0�gW4��*�4X���}G�T�&H�D؋�D�ģ�m�k��z�����Z��`q3��G���ڪ�Ɩ��Sꕖ�w�4��/G;��d��x,w#���σ����Q�c�����n�	
j��b�ű&�Wa=�]�L�K�iſ��XP���F���1\�d�����6�E���}�@�<K�u�Ä�A��
�JO&~q��[/��@o���!DXt_ВC�o����3��~K��T�l'N����}��u�ϫҽ�3Z���IT���7���E�ο֣��y��	�ah��x��l���x�J\jP~���G(�B~=�?�-�av�ba�"?�m>��%j_,���(�/>��3aaT����jqiŴX*�	U�r��R�OL��
���Ʌ�u���o?J�K���p�
��-Elr�#���c��Abr!-�V�K���,	� 3V��yb�O�]q�)_I�^�f��#��N��469��T�ڙP�C��*/�׾eU^|��%*V�[���-���IQ��dl$_��2���2^�_��z.\pKJv��K�.�˞/��'/���K'"#��M��U1��|og���利��d��A�j��ycP)x�V�ŗ�l@�٠�mN���	9��f&�c�GxH��K�k7��EJ��^=�,:W���@c���]�bPd�����~S�~�b�R��#�Vd����Fj ��?�>3�Pu"~
e	�y�/F/��ӿ\w��
�v
<"L�L~h�_���_�}a�|���8�d\���������0�/e|��?_̞���KuR�*��2�C�u��v���k��\y���~��mz�P\�?��|����7�\BT��vy�������0��YF�fT�I�oh�#��ޥ����*�8��ݧ뀴�h��`*n�W �y��f��:�(��ό��>QEv���X�����=�U|Ӗ!��׌��+63T6���u+wx�i������
�'����u�]!�Tv�ؚ��������E��~��6��~a|O�$�8mx#`�j�݉�� F^~g�c �_
~���/�闈Lԃ�_"�.�X���Ӡꑃ����(s���,c4�HH�|am�?�׀e��'^��O�'�+��m�!�nv��5��
Ϲ��㍓�M��+�j3��'�	���m�1�c��sV��r�P'틽-��P�O�d]�4^`M��� r;f�;�$���lR��<��m�b`���&��Uz��!�ecg(N�~U&Q�.,"@Y�s��#+��h8x�ֿ)���Fկ?�o3f��[���܏�l���^������nU��o9R 5��'�'5_Z#q��eY8�۵��CP�o�~Z�K���������$�»���L�NQ�dݴ/��`�1�Y�<�09�m�#���0��W\Hd�dG����G�2_�,ñ5Zb**���� ���P�Sy�"-Y��k�i̠k	�I)�幹o�|n7wr�@>��=0��������w��n�c@���/�D�	I�0��P-źx.7츤�O&��	
�r[��+��{�	��0Pd���,g��[�?����/�����UM`27"�-�!���?>q��k�FU�%����j����]ẕB��/ .���X�S��NC7���0���>x�6��O��go��$Y�{��f�U��^�ZZ:UJ���7F���o��8#jU�����o�)�+���,o�y�(�n�z9Ddb�9�zcT�
���lA����r>;rV0��S-Q~��`� �v��{�ض�F"@��W���=M-�!U��bp邷`[I�F#�r�N��G����6L�(O�|���ILܰ�dE%	�-{�]������Z��f�u��
VF��@����d��)x�Ė&!'�V=EA�]�U����ڔ�I}��S g"�	�@y�HgB�tW��#{����eä,��5R*ǻO�7Qo*�������ط�g�_ "zJ�n~��8��V�|�2d~�R��T�:�i�7)E,���ϒՐn˶��L� ]{%ҷ�ho��<M�o��mQ|+EƸ��?2qA$AA��F�RfO��@vڵRZ����ߑ��`�������H+59�ESi��f�� �>�A�r��9��VB��CˊsZ���ʇZʑ����/��~���x	\D:�5����^!��
�d�tXY��W �Jr�U�F�Do����yK�H��'��];���Z)�C�P�t ����k1h��R�iBy��# e^��8�G����*��O���Jak���,��<�"H=��P&;(eW��d?�ԥ��8]��wS�RyF",l����?������ �r�pc)ˮe�S�b�J���%`(9kN�ԗ���I�,����"���
@3�7���߮]�m�ۆ3�C$7h$ۻĢ<6�q�ޢ�%��$}�{�t�3�RnrGN�U|x��;۝�����%�%�h���N���Sb�N�{B�p���I��E$;��ǲ��En��_ܻ3��
^����#�^ ;�.�u/���֋����S�c�s�)�� ��
1Cw�m���T�~C��X��}���<�1G���D�/���?�<0��;�*���V���ӟ1���^7��=-5;J��s*k�1���0����ф�q`���G��S�a��oN�׹���S
���S**�q��ǫT;��W���JK>��|R�}���%��ha]����aUc5�~L� �C�G�d�L��.][�ZG�3M_�.6���-Һ��6�����2Y�&cQ(�Uu�*#�i����FB�mޯ�pA�xXb-�����5��+~9�o�=�� U}�J�J��F�Ѽ�#���ܾ��i�˴��;�A����7]���a��zwFj��~cd�*��^�yd^�������v�.;PY�PY�hs*�&��;��hѻ��+~{�yRK�`���T�� $���0���N�u�O�'�L��Y��ad�M�����c���Bk���S�CC����h������S�h?U�b+�7<	���PfIe����w����wn��e���x�ɫv�z��)3^��F�r�ׂ��Hz�ie��O�_�w9�}�ʉ^S��/P�ډ�q7���A����7����%"l�u�L��F�o%�٠��HW���ƻ������뛫�c�s '����>9�w�m��I�ʤQ�"ыwl�h�ZD�*��jgF�s�!��HoT�%C콑dN�˲�Άv,��yq���?�*G�˙�R��g��
�0rļvX�߿�/���������gO�a�lcX���|i���OA�},��!��?5��Cf�IS�0<z*��]�&z0�醻�Ķi����K� ����[�n�:|�y%�Gը���5��K�LM띶�t"�?�F���P�~S�{
���U�A��dю����@[��C�z��ZϮ �B�!O�y����N3$��)*�'������>ʴ�qv�^sob��f�i{��%~��|�.E��ՆN��-���;s��?��h�%�6�W�!���g��X�F�FѻDmB�c7O3��:��4��~<���a�Гͫ�ȵ�k޹SS3`U<z�]y&PQ��A'^�U�ձ��φC���ۤ!��r� c`F߾��"�u
Zg-�bK���<�6���V����ǏѢ;���	�vb�ɕ?�����-�ۙ6zk��l洶VK_��߄�f� ���W��]BWbG~R�eP�'O>�ݙ�XJ�5���3���fW5��r�{�����1���G��������#����φ{����A���3�V�l���zg����P�-p\-y	��p������W��~Q
���@ӄ�"�`S��_}p0i�z��%Fɲ�+��Q�����nr���2?1Mx�r
� }W���n���ycx��Dم=���"�g���%0��9l#7J��x���嵌�|qY�C�4J U�TyC�\��T�
mL���4a�%挟�p���b&o��7��[~��3Mo���y<|��I�b	�ҁR�3�5����`ե����~ҎY�?��u#�\�f��d��qp�
(6h���b�K�/W޲��D���<�c�Q@Z� ��(X;uׅ㑬Os�",�n�a�������9�L�L����7T
y--�^_>Pl�L�b����ɥ��d��-���g�w4�0v��0�z��e���}�$��o+�d�e���3�,E&(�](G�NЁ��P#r�Mi�YN�������}.��V���tw���2(�6(��O���v�V�R��FRo*�b�d�� -�Ρ{ �q�=���7���l�;�9�O���M����*t.�*���,�a��U�!,Nd�vd��_�4bn��'�U�{������<�^/�Ǟv��|_�{��Ӳ�3B�=��H,�хcЄV)xk}|P�-�O��6��LQ������f��ň��@��& ���9��,�W �#��dMQ���B?rI6ع#jB%���&՗��w���0(��-��Jl����=Ίl��4~U�f��\ꡥ�m/���-�U��u�8{L�`t�I�
?��$�z
�t������!x�l�l�A���b�Dz�:sʵ��WF!��&�Tm&�cV&5���R� ��i�d�1a p�sE�[60�DEN߁�P����p���T-y�:��N]V���_&��7��P������ oE�&�0�2�J��^�}p�����ӵ�Y��h�b���u'�l/�7�3�A���B@�A�*�����z��uHZf		��u}��ߜ��v�?�f�H���Pδ���{��A�~,�E��>?����L�|ϗ]�"
#~Aqӹ~��"���_�
�o�qӊ�5}��Q����{�"�3ɛHBZI�҉wj��I-d�;c�?u\e6-�''��ަ`��m&F��π���^�Л�[d���#��[{�ܯŗ�[���ɳ�H�Ьψ���g��F�W����W�&'^��&c�`�e�~]�'yH�ۂ���b���K�n='`d�n]�h�E�Du*nLЙpc9괽�Ʉ9
�V	���Ϟ�ѕ��W3�#M�P�+�~h�1�C3��.]-~/��F�5V)̥$��b��`����Sl��qskȷw��z�J�}+��*����=���w���Ar��@Z�a�ֱ���{ս��1l::�r���H�D25�?�#��?!k��si7�zǶ'#\�Mt�,��A�e�1����k!�~\�7o�X",<c��$�ntz��NLy���s%g%
XH+^�p X^�ya���xh;h�}S�����lktv�ئ�J��P��L�}�[g�uy��X��v�F�4�r���g��ڱ��QB���������'���	6�xq�����q��
�mS�:E�{	6����;��y�h���!�����d"�c��NW��,��f���^���孁�QQ��Z�e�EQ�:".��$B�4z��z� �]���X�o���f �A���0�q�z~��-��:˂�r�)h�h^7g��^��{����Nb�I���Iq`�RG#������y��J3m�U~]�L��]-}T��me.L���Z������J��D�R�F�v���~�ٮ޷s��Xi7���ڐo�+��s���0��p����^�0yz?�S�
iD�8.?��шy>8���Ip,�ڳ(乷a�b6����1��'R�0iW�G۫�پq�F[�0�0��.l���-Ti���@$~�U�| x��,�G��g�\͇��G��#GJ�K��)�!T�f��4{F`3뽱Y�l�c�z�&����oa��h�7��b|����
���E��ju�+���ل�Џ�cd���C�_ m�=n��Υ��8/�����K�J X>P������㢚��\a����ߠ�y���rk��n%/^sz�}�_���M�C]����kT��K�n�cE������0����d����K����a$%r;��c1�h�
���*b���`���/�t�'m��[ِ>�,�ɽ$L��f���(�7mr}[��1�L�}������\ȫ��f3(#���2�jH*Rfmg�X8}$��A$g�{� ~�0�8�-�$��������O�lR*�$b�g���#���Lc'�V�T:��yY���m6)�"�Q�f��I�IU>'�ɖ3F�x(��w�N��Z�s|`����)���R��A�wu>����Rh����	�rN�rn��?(d�$d�B�+-4���#�J�0r_d��Vl��Ϗ��:q�Y�= ���Q`��Vl{w���Gj��1����~�+9�;_�����l������H7�HwJ���)ݍ���)�-9t�]CJ�J0���S�����9{��Z�����yl�+����5-?���f�������o�gޑ\t}_�o�|�Z�¦)�4�
P>���?�Z4��9~5�4^TD/�ٌ���r��py�pX��u��U���L�����2l�/�gח�fO]w��Ν1�Q�/�צQD�^<p�xH��4���;J�����W v�7��������<��r���AlQ3{y�_-�9	ň�,"bv����P�a�T���i@�	 qF��}|�B�[�5��⋸ú�������Y�]��ջ�Z�Է1rfk����|P|�)v�F�uGWĝ�OI:�sβT� ��'�8����a�GQ�h�h
M�NR�/���,kc]Fu���)y��}
Ox��v���.
=;��J�ٴ'��2_gYr�U>�����ώ8���Ыw�$�89!��@�\P�o�W7�Z���� ���⎫����y��nM�MVz{ �#:��逍?]Xp�f����}B� �v��IQnt{*�c�P�6�̋�`p���/�9�|�*�<���$������b�����+`B��� *P�a	'#+	��Cվ���%���
W dm��4b�G\<X�� Q��4t��x����)��"��)��qӶk�趗O��iC>dȦ�a���ؐ0�[[s^#5 %V�����N+�=�	u|����[��Dj{hI���l�?���˼[�o�QE�(zv��u�V�W'!ڤ؆�Ł��#"�z�_�����x ����nH-��t��,�G@m5݌�&
B��� �>Q�ۣ���K� ^�4=�~��`�J��Ugr2��|~��s��<��{�Oݑ����!���o�?�L�&[���z%�c����D[�A���O�TL(�\~K)�} ��Fk �r~S%�*Q�JZ��(y���=�L��$�j��, ���3�=P�;�"՘F(a��a�G�f��7A빁�b8ȉo&Y����8��|5�	ScXaꃸE։	�AL�A��	���-i{+�������]g�]�e��(�s�։b�0��� =�f��T�jB��V���^0���S��G:�ĖQ��ՠ�:-��n�*:����%��f�؂���瀎[6�/��H�j����Z���e�+����3��7�'�%~U���"D�S�#8�R����7��G�h���ҭ�~Dч=!@q�pC��o~�4
��X�V}�~k�[2T�}�W�Z� �oMY���~Hk.��p�$�nA�`K�R\1��dZ�@A9��FW�� �����ۅ�t5��(����d��:�a>9�r����z��Aa�[-5�6� �߈��)*p�M�,�7}?^9�u+���/�JY�^���#6d�1ˑo��\�a��5�Qx������l&�XL�%�,�@��,�7��8Q����=e���Jɥx���˫w��ҁ}N�}b��0�RL�sKI-\\�YV'�C�ȵ��t!�W'���+s�B�-]8���E鷟QZ>�u����#��G>T���%��W��_��S$0��-�7Ok?�FY��|�/��z�
��,���|h�q2䶐*����$�b�^7��D��(m����&^�A��)�%s�x��y�yͦ��Ș���E�0�����9Y���_�r���K�D|&�1�w�Qz�X����2�Ai�B�Jt[+r�12�DM	��燺SGBxtf��oQ0L�"Q&0M���ְ+D�S�v�፾��� �E{p����B98Ȓ��Q5�*U+Iv{�s��U˒�����`��!v�k<����-t������f����?.�;���N�&� �r�T�!s�	輶�һ�P�����#_���:�_YZ�X��ޥU<A�s����e��\)�6��L�^Y���D*P�ڴά�Gޣ�9���O�]�l@�a�9@0�ڟ��]ۈ����R����i��xYO��Lk���o���0���n�	������Q�r�n-v����z�9��cB����-��ڏ9,�{�)$S�S����\.%���$ �CG�	�?w�2"}b*4�
 �d��K�����-��k���T}���� O��d�0�_�8���b�>y������2�[x����'7�l�e[<����-�h��G~�Q��M�iԆ��h	��տhP�����@`VT�y�}�[l�y/,f�D]�
�==Q�i�$��l��Ե���^0$�,��[�e$mU�!̻��� 2�����L;�5�ɆfٖkK����📂66Y$��O5��O�>��9k�����r[Q�l3���D/�[�u5�U��Ώ��xf���9�<K��ϕ�:7u�b��' RC*=�O�᳟�N�D�G*�鮀�W� ���p�v�A�ɘ�_���R�M���jԚf��.���I=bi�PvP
��rf@;�G��x������Ŀ0h�gg�?h��0����$�ɉB��+�u,E<�#����d�W�k�቎�?d�G$��`��Se>6Æ)��'���1Euv>�I4��+@U���Ji98H��:�,�n�p����P[�h���T�=T1sżGe���hCȘ�N�af��������������l*Z�������_t,�m�tA�p�Cא\�>����sW�6�ڥVb��%�ĸ�3��&>ͅ�p�va��?���[��2�}�J�ɟe�cpP[��!&�n+���N�1'pd�w}�����
�O>AU��HM��5�!�vU��7�	QӠ���RI]��ג�y�ۨ�W�St1�m�=�At/��sr�B�_%
Zr@sz��^������ �P�vSǋ��eI`�WY�Y��+`�!�=��|���]�g�7�H����*hٯ;&� w��9��X�;��Ғ�9I��2��;[�j��9{��Nc��Tq���)�����h�٭V����
5F��%�A��.X���^=�}U��0h ���*�Zy�l���ց�ٖ��fB��)H�P���QF�m3����E�Z�`�M����� N1�M[�ʽ��r�tI t9�:M�����8� ��u��w����;9W��K���u&�c�P
��Wj�a�;�W�e�Kb�צ�[i�/�b��$�Öe�x �SG�i���W�F�Fލxը�K�Iݐ�&������
]�Nk���	�[U+=�
�w��f�`O��E������V�CT�_�"�� W���>�&�NP.�n@ఒ�6���y��Q?�޷ӹ��ZŦ�'���(T]��c�Ҍm�o��� �/�[lץ�����t�?g@��途U�܏��%u���꼠��)����%���D �\�1z3H��D|�;� ���
]�b�Zr:��}MU%8�H�|B�7�����V������U2��uL�=�$�[3/��?�dA��U�}�Oz�����'�?��vm
�}s4G
b�o�$խ�������YaP��5X�>49���S�L]�NCA������:�1D��������wU�/�����q�)I� �|��>Y�J��[��֩�;�W�QRퟆ�P��c)������q����G�\\\���7��C��®�A3J�|���7@�o��Ѹ���H�"�C(��ڐ3��*� Y�B��q����z�&�F����8�cQ�G�����S>jk��}U�H%��S����o��L�/�N�{X.9Q�R��̝۹�y͏ܔ.:�EƲ��2���v~��/��Jʝ�
.�;͔~(���{B#��o�o�b#���3��1��Яh�T����g����rB��]s�,T,��-.w�n"d	��Ն�:`\�_�̷��G���K�ޟ!��� ��>�k0L$��b�ͷ
ˠ��=U������qZ�bt��{d�Ć���'���Wx��C��qĵ����-K��Ϙ�oR �b+�o��솉)#����kITz�(r�~�@�R�O�k��y�����B��T��q�ᣫ�Խ��5��i7�Ku��jB�UxC��-����B���``l�`4�(��<���Vؐ"H��YsôehNS(�w�Q�qE���2-o��8����~l�7���'?A� F���c+O�&���3W|Ց�ld5���B���ɘ-��M�$�1��ڞQ�8�C��n� Ѓ�� � �ɤEޜ����1E�ܫ��L�I�w�H��Bg����+�"+���*@g7�,���˵}X�����SB�c��)2���/����T�{B�v�8I!��%z�/�1jp)����Ʈ�;�lx�5&מWݙ��㾺�92�x꿓�����[]ڰ�<���7_�N�$`����P�[]u�Z��@�<>�v�s��P�����t��CX���}_�wi�������*jL��L�������
{�Í�prY��MnS�DE̻ٝ����#�r]L�W��H�No���$���m�K�|�x:�E�}�5|�{�<)bś�����g����W@$e���A����&�9�t!�����鱁��ˎ��n�u�����ٗ>{r9:����)������+�7��z��)Ȣ�-/?�u}uc��=Ψ��4t�~��~�m�}d~4g3I��9{�ܿZ	*�{�:?�ְ�1�Eh�������]%��^6�t��B�>k���{<J�t�v�;�9�P��޾H��ynj~�:�]6e��S���Q;��Ȗ��N�]?�x'3v��6���gD�L��X�mL���Y���%�u%��w�ƶ��j��I��8�/��i�gC�/g_u��o����d�δ%�n�*%�VSR[�@���*�qx��Oe����~�������� �vmrꎌ��I(n�����	1��Yb�ɾOѳȟv����kT���u[jM�;��m�8�y�zt���p�tj��j�N�ʳb�4�����acC�.+wN.�XB�����pr;��y�~����R�H�3�+�+�p�{���~L�:��t�c�]�:���[@<�!���\os��4ōW:�r��.�X>Yº��ΕIE�*�2��K� Q��"Y}PY�^KKK.����\�{P�,��܋���Q�Ѣ�quS�n��.]`����}r��=f��A��S���Q���+�VL�"�m��3�]z��>����~��Z6�F�������έ�yݝ�����gEwؑ�8�R�*��Q���p\��PQKj%��ۂ��<zr���c,'c�ɟ'�y�؆�̔�["���Mkg�k���?�R�y�\Tq��6�2�����h��Mp��V�l�ƅ��Z���~$�|`F��4l�?Ğ���p'NkPDB����|	��kst;UX��ø0ם*����o�ԫ��������B�n��l(	����%�
O���f_�y&�=�*?x�
�M�T��R�@� ����9��Φ�c'��*f��d�g�̿!��KPtB��=��p���JcC<ڿ�����lCF�s���{/f�ڎ���	�\�(�e���h�ᇍ^i�XT6
*��-a���D����z+���p��H��O>C�G�X�9H�}��v�Oi�b��1b׶�`�����{I>����Ębv������~P�ۗKC�����T��9�⩲�a�긳֤
�g��>pW1
��O;`t���j0�Ʀ^������R6>�G��έ�fO���d
S��Xg��L׻59V���
9�i-�O����ͻe�X]d���NT�uQT�^dk"�#
����L����:{
ށ,Y�i�k�?~A�	�Q�"�)��TYRF�(Nm�dX�!N��RsgS�D�>6>��c,��̆'�3	�������,%���B�1�I��F%���l��+:�-j� ��*gU"�
����:P��F�Ưx�[��Y�w��-1n���!�#�"�*�1֐]A���'j��P�4�S���G[#�
c��{�8�\C���_�����4���DI��q�裸E����'�]����.����|s���-o�	��(���^�{�����m�)z��W ���sG�S'�@�W?"�Eg��_�YĺY�e�x�Cx"�D�� >v{&5����(�\i��Ӈk�,�{��]�ApwD�a���״}��M��
���	�iY?��3t�$�����5��/Xs]�@����������t<7�ݥI�o]�m�AG5*�p�K���nT�)>��(n��+ Tr��Z�FU�Q[[;��C�}J�U?�Ôu���N�4�Q�8b���%g�����7���-�(\䊾�m�H[���r��ƞ/�5�yf7r#�%���wAj^�Q�،4�@�ѫ�����i0Y�8��0�|�	�Tٿ�V�G�p+ݰ�iR���*�ޒ�8��&Ԡ�Kڅ�?=sDz���x>�\R�"�]��f}�^1e�)��	���TV�։�u�k�Ǎ񆜚�|m��e��������7�}L��*�V�I¹�B�����U����?�T.
e�h7�绪��76뢮i73%�.���Am }BY�����I4I!�Nޢ��H���r����!R���|.eI�ǆ.�y2d�?�$55X5�	��d�%Ǚ7}���k*��&�uJ�뛂��#;#Y)�Y�W �#]�la��|mm���b
#u�L��'���ө�����l��ۚAs��vs��a�Å�q����͂\U)���ޞ��j��Ma��/l�J�������Au�_�
�G�c��\���9��d0�����d���4ռ�R��d#�cC��"����/�G]����T�?������ED�O���_@���vוPI�|O��� m�XD2�>���s��qBu�4`��p������s6��EP�7�D�Ie�R��N$��L$�V����cus��W�\��fv<���ᶂq-��uڠ��Uk��>6��Ɨ��?����،����;���T& L*��TҔ@�߇/�Fy-?F��,��`����5��lk|!�o���݅��s��u
�V��Hm�-G��b� >��
\�v���ʃ�ѱ��[�;9��Vh�B$����Ri%7�f������og%�y/95�H��l�,��t����48����Yt>�a,�N��;��bZ�����w��:w)g�7��)X2g*�yb��8��~�Vޝ:N��q�ɋ�j�۶`�m�O���n3]��V��x���$�@ UII=���|~Hʤ�ؐs��Z6��d�L]\�`3|T�/��ۄ	���İl�����.i(*�W�|����4U)"/ ϻ�5o
�*��� ��󍒍��O}v��9ӣĢ[ �f׸��N�4�,�w]J�v<W��S����K�~���G��N3Zl�+,K-��4Q�'��p�q���Y�'�J�'@���ߓ6��2t��l��nQSf:EY��ʾ(�뾤���ٞWe?�6��B���]�;V�&�Q~0�����>�e]W�Ĵ��<P�|�v��a��y7��dD�]���_E�cȪ���h�`/�p���mr��|�����=�o�9.�ʲM����d恔!�� ^�����u�=M�h$󸛪�黔��nQh��z��R�񿔒�R�� ���\����f�!B2ȪU2�m�~�?kC��:;Z��Ta�@ ?}����M�X��(�t���c�$e���*��yR��T)M�>����8Z� 7פ��{b~L�Xv�+�	��I�:x.�ܞԴ��D@� P�e O��o1T =�8�����R�%YN����-c�Ë���W_A��/Ӈsi+vTw(?R'nFħ���~�.�i����������h����J���U�N�(����=�Y-�S��j�����r��x��^�yn���y��2l�۝�}��s�b7WH�Ӫu6?���-�BX�h�ƢX�����L��z$	NU=��6
4ڷ�t�\�aJ�<�UU#d��˕sͼ��s�ql�K��������Y0�X��[�+�W�@gJ^Nz��
�i�;0@5�c�A��]��ZE�Bd���p��L^I�h��ME;��z��?�V��h\G�::f�D�63�,��g������7��4W
�P�N�;R|齸3�\Rқi�$P����'p^�ɔ|�t��#2Mb�?�
���'x԰%&+%I�9�O�e�������Ǚ���_�>�ة����֯R���ASra/T]��D����7�M-�%Ub`��]z���|��y�d�5"���K�%���J��|�=${�q�{��x|��8\P/�H��8:�!�����R�����J��
��m��U#��!�h%J´޹:{xnT���D�n�ϒ�Ӿ������(�z/��-\��׬.��*4@[~`�X)h��|��*���~�o\��
�i�C���Ll�wƸv#��" �$Ar��>7�
�Y��4�O!�a��=�KNS�F�F'��(������Z��,�cx�_X�خ����	�H~�D���S��h��8#��(L�Y[rs��y�CU��GeW�	р]��;���o��~�8���Q֫)�X{,"H+�#{(`Q��)�_~��o�ܬ��޾���D%;����p1�^$_<N~/��S7y���r�n�Ît��d�}��x��t

�1�G�UkCnv��n��A'������-�uf*��W�eMǕ{���5?_��%�wm��s�{�7�J�uaa	�/��7t�����9��@3�X�M���dH�wP�i�[�I>����.�9]R�a������J��Vq��
��)]����_���9�e�S�Swg��_�:�<:]��s�"_��g�3'��lÇQ�6�	D����6��U~�I�"��������f�1Ers^�;]�o�7�ԅL�;�Da��QQ�rUn|���|�著۫�_�ռ��O;�diEnM�:���ƘE<��yn�N��{=�m��NQ�;3����mKA�+��'@琻�H�J��E�W�l������a�S�z��!�����(j|ބrߏ�n7����L��0ӯ��� ���p��)2U�:�7�^�HjoG�M���Y?{[�
�2�5�"M!�W��.��9�m	����������̆V����U�}��<�'�C3~DT|-��?�/(�ALA� �Ix�`��������T�q��1wkcj�>W�M�i	�3�{KC��7>���O��D!@�_N�������Ee�s/��N�w���?'�1D��=�f�k���JE+��Tco4)��%e�p��:�x�$Z�XE�uP|X9j��`��1��VU?uW	E	�p�<ö��Oǵَ�|�c-����T�@�_=�+x��Wm�X:�agT�Ge�ay���xVY�Eu7�4�C$����.ʒ�qvk2�&(4�Yh	^��7��%���-���&)fTHX�q�@�eaObL�z��!j��2�Kh�|&DStX���#��>d����)q��=��c���i�W�/-�x;=�h����><9D�=�HIU��?O�5Ղmp_d\�#��z���Q5�P��|\j���Y�)�L�E9\^�%f�"I~߻*d͎�$lE����ﾎT[�����?PqV?U�r��]�ړ��8["�Bn�{;N����̷]o��/	�Ev��v$���T;�R�V�d|%��M��d�F)}c�R|�<��O��]��ʥ�t����0���� �h�bR���Չ��b�e�U#��I>��t��B�2���o&105�mq.N��O_s�ځ�/��^Nh`趓de�7ZiS~�Q���"���iT�q-/�|I���1�|-3x﨣�n�57��vB�"V�zp�\�V���{������׸�aϯ���c�%��Ԗs��m����R��N(#���)�b�`+V�a��|_!!�EL䦒�D�&
��#$��#�X�_��U���8����6QÓ'�[9::�
�hkx7�/�+LV*��ޟ5�D�p|�6oP����E����?��ۦ��)�r7�٭�G���7�u���%���)%�*���a�l�ؚ���b	��P��0�I���c��C���qk�V]g4`�v����
�߰?�J��;r׺h�Aa��u]�iZ�����6�>��I�e��;���7"d�N�p?
��*���8$��(�n���O��h#��Y���H
ל����!��	>��5R��V�舐EtR�=�3�a&�<1�Ƚh�%r8E���1K�
�}�C��&ǂ9���񷭮s�j���c4 ����ɢ�R�y����#��� �zM�6G}u���|_{�!��z�2=l�,f�ݭ��#�GUe����R�o�J�Y�����ƬNEy�:�{G�2��)�Yr���+]?��3�^�G��M��*wVb���U�U{��،4�iא��`/)���܋O�zW�B�h�E��W�>�{�^�s�կ�)fT��v�����F���@�����s�V���jH�f��i��O��>۴A�W�;�x���E9j�B���b�Q崢�˔>ޅJBYh�&-�^�0q�a'��,�e�x�ML`
��ئ�\��3pH�e�pG~���`{�����0�����:1d�
#��D������3F̺��cdỊ���c~S��l� �F��'�o�����mD�:Ǩ�ÄFj���w���ݷ����wSR/�����weJ���7|�UK1�=f�_`g��-̹r�0X�m�W3�Y�ײYC����S�R�-�Owif�_��H��{QrU\a�?��ew��ފ��1��J���}0�'(�A?�/�ݍs���]K+T�d��tѠ�Y�G�V���ӧ#S����C��xn��7N�޷,��\�Lf��K��͝�f;�<uDݮ���|XG�+�n�u�f{e��[���$�)�S�J ��Z絾�fb&��]�~��u�.����Mƈ���Q���e<��ef!��)
�q���o-���L��|Ntؔ��� �/MY�-B	��A���K`!�e6x�I�T֡
��\�@H�N��L8�$�5,��l]�E��Rs��[���3&��о6�f~o������Z�=��z�~qC�95Z��:6K��1�E��4k��deRq��m�e�XC����g��7a��_����v�:�I~�r1�#)>��
�=�u�ب�����i5g0� �-9P��
�
�ǕCl+澓�cw�+$f��0��.M��  |�P�V��+��?��'�����Vs(�]��M�0eh/��4,����$K[T���R���/-<�I_�E��J�S��3�Ħۦ�����HL���U"��d�_��ר������[ˁ�m��B-qi.39�]n�%������:},!!8���8�@��:ٖ���5�;U�i��C��g�
�K�/��+���|��!�r0i�&[�9�^��1#�a��+;��رIE�[�j
y%�{*��6�?,�`:���ߣ�{�0Il���W�d��4ZV�c�Un;�"=�\����^%�Х�*-_ʲ\�\���Ћ-�!�9#�������b�z��Yb#��_ՆW�{�Pk^a#qe�Һnmʹ6��O���uB��xF-��f�x��	���<z���=ۗ�	�o#��c���!�� F7Q��U�]�����P�
׭�og���8��H��Ǘd
�k7e��_R��b*���TW�Il�]���$�n&m��b؊T<����i�T6!��s\���� �P��������l6;�w��j]c{���9Q��W}UT���Bηol2��(��`*k�񡀹��W@tb������;��,A��~��� �uf�ݤ�"ՠ�mo��c5tC��m>8i�xx��Y%w� ���m�Pf�W�:y�Ó���8���|�̤̎Qf����M%O��x�A�# t ��]���R����A�Ӕ����n:\4�,i;6��0�zL�"�l��r}h)̯6,~6�.��CgLq�T{b��6Fy�c�G:��2\x;Q
1!�M�2�3�3 �r��L~�����\�  �ػfC�^� {�N�D�Z.=���Gz�ur��M��4d�"X#L��0R�^\�y��}�����wu��W*=ן]�i8 Wn�g�j�z#��X�2R2�c?��)��.��`ꖤ�Wi,ˎ����p��j�<�=h���<�P:=�0@˼xp�����ؘ��v�1����_c����۟+J���[×��)r��/p�2S1|фI	;\���3/ah�>�5	�v�`=����[��2`�Í���e�p��g������21m?��@��j')�� �l:?�x�dxb��{�2�ۢ�D&
n���]?�x���߫��Y��=�PM]w�w�Lb{�[9��V��ѣR�ԋ��88�az�y^�����k&�6��Y���H��0"�O*b�{u�%�c���uʼ�Ө���lf�<��X��Tům��	_>�� �����{,���-'|��)?{� w�&8�p��o��&�����?H�="���*��\��Z|��}���d�1n'�u=�_oQ��`�|DS��..���v��d�e���{Uf��g��ĳ�Di�;
�'i%1��b��-r���ox��+��λ�,�Rg�#�U%`Zk��_�{��FH^�x	:}�6��t2�lĵ�X�7w6"�R��3�é��cS�Œ&^i��h*dgs3yE����J�G�0�~U�41��8�U�3��j�	���@v��77v	������}&Vn��H�,��V�K}��l5@�7	�Y[ht��� �[��'���)���R��%�"a�W@+,ÊXF�Dw:�et(R�>5V>���0�|V�(�N|֓���J�e ��6m��+�铱Y�7M����x�K&ֈ�.�Λy�B�1�R�|����F{�`\�����;��Y�#�W�p@o��,@�4�9f�r$Oe� �wTO�.��*n@w1�cj=�?Q�SߧW�O��P�q�e,���zf��n���P�����b��7�qiL����{��]�0MS�_�sxyu(V�տ�	�h�*L<�D7����� oa/!&�v'����;�����q��(N.b�_��]<�6{A;-~�[^R�����/��\i�0�n�C�uy2$[ŰP7��k_��:l�%���6O'Ʈt�w�k�Ƃ�����vxY8�8j�U��?kC��Ia4�>߾�l�U�����1��U��Ge8Bi���Y��#�	�����ġiD��վ`���c�0��h��/[�sTY��hXm��u��Cz{����d>�����@x6~ʮ2�	s��3��x�Q1�Q+���c[5����mq߱��&�q#�Xz��0F\���5�����
,�`�M/ZY��f��s��`P��ڲ�	�nQe!��Ì�SwgƗ�����ȉ��T��Y�����,��j��_�f��tS���*�f�(��e�}���v�-��������:��� �B�����M%��B:��h}ǥK=�K��A�}��=�����!����tv�>��W�v,����y���ʑ������Z��8湸<�{Q=�xR
X�Y|�l�6�ti�a�w�_�Ma��wt�jYɢqѢ���՞k�@N>g?���K	6Cy��f�G{1���t�%��2ܥ���B#��Js(8��_0I�"=:�q0\Z�F��
����&���W:|9�*����Y�[!ȳ+1��ԐG�gF�נ\i\�j�ي�F����>D[�@���'�����#x�Om�%��d�R%�˵�CO>�	�y꒲DN8s�K�+�˸���%����� 0�1�+����Jl::0J6�$�M*�P����({�2|�ܛ׫����V�Ce�'�i�Y�0H�"�%%MCYE>���*�����V�g�_����W8�:L/Vn���|ɤ����I�W�J�&��{�IC��TO�5Ǡ3t���Vn��+�S�9�~!ٺn���j��V������6jܢ��Ǡ:g�.7�7� =���t�h���hε�FI��Th��*2n�ʷ��6�?X��*����cɗ@�����7����B�Q�X^Fk�5�q1ԭU��������eJ\8�n���Ae���K��u��7&%�v�5]��%�K/6@P��T}=&�/o�2�Բ�p�-$f*���TA��"�����a��ܤi�O8�b}:G2���oL����ǲSD���G�e<��p��*�֩�Q�u��~< ������7D<��x�[���F��j8�	4�D�^�
�� <}�"��ҐΉ��R7���`VE�=�KG�S�V ���a��.��{���J�%�+sr�&ƹ<�]��h�ЪGq�W�cMR�q+��3[�^��>)�6G&��������G4����^};E��N�h�E�>�zr��sB�'����oӼ�s�Ya�[r\.��ݥ�y�Sg�RPU�C�n�4O����h��`)�]A�r�i��>4ʕ5�Ҧ��rEk��s����ApK�5#X[o�/���?�#�w�ъ���i
_HnqUm�/�������)��"�<���;���WG��%���
?�g����K�$~���F���%В
���z,Iwu5��\�F�%��#݃���������Z���W�ÂI�!j�� �䠺�U4�Ek �Ǳ����5�F�K|eG����C��b��a/�q��sHzޞ����;~��~�BR�H�aY���
�yi�)f��~�?;��	`ӣr��#�Np�Q	�9ӫ�eƮ>�1PHϾ�qB�BS�{���L���6 ��g܏�<����4�q0��}l�� H�X��R(�c3s7�ę�v��}Ħ�-��KFl�Yl/�=�iʋ���dJ���l8�n��LR�Z;M".?k;�u}Bp�c�.�)CP,����1P�;à�_�I�
eJM�oǇ?��чZ~�'@gP��8�a7A6�r�:.�MF�2򑮈�ކ�s�5̘vt���#��x�I�����"���	�V}|��OB* ��D�[=8_��IU�����m{�(2��[_�/'MM�=��yk�SW%��C�M�L��g�!7�7�W-`״���׈�����&rg��U��J�����h<�1�%�Pv��*�= )�j�L�w4uy^�D�|q��
���jY)�o��&��-̈��G�(���gX�IQϯ�U)0��oa�:�6�+���ΈG�	1?sٔ��a1�zEM��mx�lT��k*X�F��?91��sɢ�N��B�/�6ZW�<Pj��zM{�C���Y..wh�[C`c\��%��+��A�c�X��J�_���Ah�S�����rQ���{e����M>�Ē�>(�m���=fa�hش���y��r��^��[�%# `ӹ^c��o�6��g�f����8�e���A�	*�O���
����q���5�cgE����;�:��7(i�/j�Z��ĝW�$O�$Y��4��pdX�n�ɺ�o����œ���I:����(c	us�T�����#�a��G����N�^؀t�h�J�x�ȧ������]f��IF;�v<r�!yZ�
$�"�ӟ$�0�_��G��7š:��#)bA�u��Lz��Q�7���D�;	׿�U�#�R9K��Xq]&-��W:��R�*��,���:+����{�19ʶ?}��飻�z��8�Q��q_�[��KQ(W������8��Nv�0$iЦ�B�@����=R�Pp�Ӗ��=�I��5.@����4�9x��x�z�����	^B���;��F����\${��}V�K>��&�Rb��>�"�N�\��7�c�<Y���D��������C1x��15�YƦ���C���ɥi?���n��d,*�I�	���]��6�#�鴄hæGAZ���ǈ�)�7�1�fh� +��Cn�VB<��mχ�NC-ei>>�,�nw�uFulQ�?�ɓ�
ޱ9��q�UA��;��^ꉛ���3�f�gF����h{���h��;����тri��4锢t+yYv�wSis�1�̛�<v~��'��Avu�<�v�'���|앒JK3qa�("��vu��+)����xcM-4VS!���h,M�� tv��!�ȏ��$�,���wWQ��z��p�/['K�han�o��,�3E)����F"*t^��kK����Ǔ�r+
�l���/i�KՄ�ӝ�>L��t\��
����L�ݩ��0o"A�������ڋ�� �u���j��.hJ�N񲸯)��s������;˦��`mB��.���mp\��www����6��C\'�[���s��]�j}ؽ��{uݫ��T:l�X)�[)�o� ���v76X$AY1�f8��~{�üu�Mhd�-����E�H(��_�߭)���δM��w�/BT��n���Κ;�	�(��Çr%���P����@��9��>K��;@&�YP~��޲���'�PpA�n<m��x��T�>�W��ҕ�/���)|�:��3"���Ռ�!�jz� ׯ#}g��-����6��Y;:5��i�H, ��S����cC�P!��<5Mi�,�4��gu��[�y�S��V��p�$v���������"��z�����H�s#�I̍��0���L����B銳&�&���p
����؍�� �e'��I4Ь�?�����v)�H�w��U�!������'�S�On)��*�+F�r�;Ȧ_f�G�m"y脲Ԣ9�e�90��qA��I�R��o��=2������,�*�?�9zf�'��s������0��An(�X|L����Ԍ��ET*�DD5-m��%�.V�&����w ��+Pwy���s!�Y��v\.����g�I<#�l��a#kWF8=�C�Tvor~�Mo�8�r���G���3sa�ψ�#��Q��0�4q��H���d����P'�f%k�`�Ho�+��*������1�\�C��c	��;i=�R�>�b�0s��Fͯa�H�	dr�D�;F�E-]a�![�
]�S����)q4;�#�S�DC�0�F�g��eq����&��e�m0��0Fs�[\����Ǘ�5w��4�PHs�OU������_�ؙhJF�b�='�J�Aɦ�ړ���#�<�]�,)K�wؔ� ޼���do0�B��;	E��������ը;ݲ��5G���:A"��1�'��Cn��{&.e�\y����$��h�TT�D�1c��#�1~�/2:熂��)�d�E��@�O�}<rG�b!�'%!ڧ�K��ج���ta4��hNyֶo�T̐��&%eoև����߱4��̥����9A�<5�&{��er�K���  GP�ά��{�=I����<��$�^�P�"?��p��Շ�5M^}l�|�0E�AXY�2�#��/�=����jVBTxw���b}ϧ�%P��Tk�q�e�᳁]	>�Gv�>x'k'�9W�?��;�#�Z���'q�J��_Qӧ�V���`f���;�ى7V1��&�e���*F�hR�����k�*c�~��nN�Y��[1�$�^�-D'�����o��5B�ı�ù5�1�~1�@5P�9��R�ʀ5�����n-��n��z���ίb��������Zr}��1���*Z!`����(��|��BӼ���s�X���¥l�{��V/jR��I�~P�~�|��ʑ��M��>|k֮�6�ۉU�%��S��2�ȓlN;$��Bv�*r�B}*�JMmOv�1s�@��?�\@�O�#��aցN%�%		�|�y՗J�rlf�Q�w<��NL�#k�at�h��S�L_��bJ;Cܲ��zt)%��p罀@�+L��\O�5���@����7C�i��-�L���'�\76����d��;&�5+�GC��
 ��61SۜHVz[��V>JQ�[�}Hp���m�&��#B?P}R/�����Y�}7JFC*/cB�)vS������)��O"�������i���㨰{��z8�Z�D�1�9�"��)�x|��))[��I.��k4�N�L��/㞓�Kh�c���PpB��m�et��K[U�6���F7��n�;��>�9D�_(��1aQ}�+�C'{�r�:]��_��V�"W�o�J�Á��դ���3r��<����z�3�}v�Z�R��f����*�k�ӫ�������rj䰰�2�򽑔�1-�.��QZ[��z;���u~O$���	�o4W��K.GͻL���Ȋ�u�$��5�]�z��NW���0F����Y��o~�/%�%v���\
�L�B<��w�C�[�0� fĤu�G9��i�?F�o2Ȯ��F����\	hF�b L��X��x������g8\��]��-����h.w��l���F���0��ӛ��V�r������%=���<���}�_L���r0��h�i��(������|�§�9�K.=_��ȓ9��fw��|&vҝ1|�|0>���ꠔe��5��L%�-\�.*3�+i�o�٪�H��%J�u��˲Wzv|�6{ɘo[1~Z��,U�
%�� �/Hy�}�%hz,l���m�����p����<�C�XE�bglɚv=���mK�/�y0'b������pN����ZL�=���B�e���ؾ�k͎d4�d�S��o���1���R�r�]n��{V��	i����&TT��N�ؿ?`��\��ɗ���v�z�i+n��=��p,���f*
L@�Z�f4�Qz�h��З��+��n]Y��T��C�c����QH�_�9;/��Q�n$�F{@i�4�X[�dXy;j��T�n��n��$���2E�c��#6�!5\&���>�{s�ܽ��q<el^�� 'Z6���oiz��t���;ӯ�l{����n?f\F��vAD^���ߖ��v��z{o�ix=e�~�D�K֠j_��\:�dr�bV}�Z�-���޴,j�_U��ҟә��V�[����+��|~}*��Z�$Ϳy��.�R��<F���v(rmT������A�В�V���x�BU^���yD��5��NR���zg}��F\��x��O�)c;�_R!���0ݜ�������F�U�/��
Ȣ@��}��[�
ҫ℃�ƚf����T��*g=TJ��`�m�8Ia��B��n~�P++d�k���W�4ٽt�C�y���?��fB���Ͳ�P�1C�F=O��X����`Iv�E��MfxhK��I��3�޶%^���&'�����v�n���5�/DO��a^D�@�5���3	�>:G)o��b���N�6�t�0����n�_^�+��g��S�!��u��xjJ�� G��g��(^<��蝂���6���ТJ~�ZF�@M�Ct+^7o�Cn��c��Zy.V�������
�xH��\l+����J����4����S�ȕ�R��UK�f[��>��Q�0�؟��㛴2�MY��i<�ک�Ȓ���Su��g�;!)����p�����u���IOwGvA��]�/�2`6�XV��*�EV�#Y��!��MFl�4r���.��}�s��܌�ο<n���}��h>��i�!ڰ����U�^�G2�;�2"ۄK��ӌ?r��jj���i�R���_�����F�J[m��k��GŬ��.���`�4�'a��7�Snr %X��n��0Mvws�wj�`�E�wm%*CD�z���~��aUُz�M��h�b)sX%�V���-�)��6��BOE_��) #CԼg��b��g��}Ҿ'�V.�>+JB�ُsog�J{����
��5Sc��G��lI�;�������Gu�4P�Yz�ѝ�zkV쥎 P�$���ie܋�OڤC���|�ښ,��ۖ�x+̮��90{�}�hy�qs�q�ݘ\��X^�ZjͰx����
xҢu��R�k���������'�e.�z[�G9��HMg�^��䡔�Q+�Jł���pT�1�Nt������^�z�rA�_6s�j{�mmj�"��O0~�����t֦����j�%�/�SًВ�F_��4j��ÄS��8�moΈOy_�*f�@��EODz,�<��ۖ=\�\f�D8Q=�S�Ĕ��K=n����d(�f�N>%?��vn�o.��$���\�_��[X�q�؅�wJ��n��]{�O`��$��Ҥ�o�.]��.^�J�CW%Պ
�.��6e.���@�a<����M����T<��I�(�e�q�*��28�����ݫf~:#�L ��E�Ip�~����� �|i�ȭ_�����/�S?:�_
�i���wm]ͥ�m�A=��"=��Ll�D칊��R�u��o ����.�Ts�^J�^{����.l
$�O��[�I�VPŽ%�Q�Ƥ;'Iu�E��T�yw�~��9��eE֗���=*�Ұʟ-���_��ۭX:w����飏Iu,�h�4��$P��)U-,����[�or����"�Z}�Rܯ�;�b�!����p@�ѱ4\�߻MW����<E$"�,�%�@���~q�����Y
�8ӵ�*�߿	��-��r)��T��ߐT��\̄�����R������2��s�v��~�ٶ�'O��㺲�Hd�V1�/���$rs��AG�3g��=�n7�I�4�S�����S��T�bG�'�pJ5 �hei/D�s�nx�-��q5�(]�߉M�{U����Ru����o~������m�nj/7S5AsgZ��୨�x����r���ʴH�``�a /]�K�%�=�1���
f�a���Ij�#Be��/5/鋉��s]�¼��56[ӥ~�]�.$�i��d��>+P�}k2(��~�����(0P�EΊ��D8�8���l��G���������kb�"�
�����	�tm_5��_@�g�TQ�$;L���Ml����t��M�5�V��y�����RA�qի�v�����(�7��dYk���	GY�HX�S�eg��Kf7&ǼFuR�^�F��NHTO�0G��]��W�mC�Ñ�y��I(v4��U��%����mB���]�W������Ib���ؖw��Ғ��l=����ם�c�2*���/��&�o�?t_�7ٺy%GمrG�[���O���ZU�zӵf� ���>6@��ĺ����O�O����n�ް���Y�Ň��z�������5��,@�ŚW���O"E��
�H7.N��LB�J7��04mM*i��4/��B�?0 G��e�w�\Y��f�' ���Pjd%>�A��T0pT���FH����|�HL�9��݃f�>���P�OM�%�_:�9��%=�<���Z��Lϩ�������w�:Z�c=TI�Kk�aa�a([z��Ĉ����4�������S5�0$p��DڮE[��)i�pim�{��Tn�~�n؜wZf�vO��S�,n���Tb��w}�]������md����)�K
.��" ~N���������M���i�Z+-㦘K9���������kܖnns��M�M�pn���׷F=���	;�@��fs��S��{��A�2��n��i�\#ȫ�ZmZr���'��6�T��m��>�8�?���] �9���p�������]����E�^
�AI��H����o�,�<�N�z��zcמ��[������>�#�y ����g/^#�f��X-�X�,���BO���l�S΃�6�a{w}�S�|sC+�\�����e�+ThC
"^��c��,� %-���]��\���:Ϻ*���/9ڽ�_F/l��5�m	��*��PO+��̋\0q�R�/]V�4]��.~(����,�C��&��/ÂZԷk�)���0d���8�r��i�0I2[�����z�j�������`�s�2���p�>޺��h���� 9���/�W���&�pO��p�ъR0�s����Ð��;�����s�u�#��������\�s�Q+s3���_!��՚�hxs��xbAݼ�;�;�B/b�M���H�;��e�P6'���y�&bϡ�E����nV^�2���rN��C�U)�2qC-0+����W��̗:�w�¦7� h��l��> �T�$��T%&k��.,^y�ק��;N������.����*�K��m��$�(?��˷��7��ͫ,���t�W��G?���Տ:�oQ@o������^<sXA;�D~{�Û[W�MOe�s�EM���C[Y�M�?��s����=��M�Z��飲�;/��������;��慠����cdG��~{�铍a�����i�y?/{�|A�IM��(��*�JET"ERH�C�H�IbF�}iFTf�	aw��.�%T2Qn�`V d�sJ�6E{}Y���Ԁ��ր�J��:��vE���2EId���2b��9{�8Ht2 9,9`pn�1\��� ��������B��A������s�6�X���h��;�����(:�.����j�M?;��PCmJg&"�H��<W0�x+�"��X/�OZx}ֳ�4���əx3��d�x����)�.�KH�:�K/�-��^��� [�`E�GS��UnH�\B�'i���)��>I�}:I�Gm�m���w���p @a�pΉ#P?�����{%aO97��CQJ�7'��HWm� tiw���7��͕���4$��c�
�g!�����ӛ��lM��x�m:$�x#ڴC
a�C�4fF����P�O����%̑�����F�n���T~��n�����L�W���3�R6,n�-��7����<!�u��,��F��I��1���̇�sh��`��*c���c,Bq>�fB}|�L��=E�f;yaG��-!��E�U湷=C�F�JI����)��sNl9�qpg3�@�k7f��	���Ǯ{��e��� K�R�UC��R��zZ��^�h[��vX�B(	5����:���zJ��v�<�����7����E�j_�O�O�|,#vKђ22[�0���Ką���|�;E��E�B�	HZ�gwG��]˅�i!Os�[�N�4O�q1�j���3h1 VT=�an�R�^��o#*�������q8�պ�*,� ���s�&�OvMc��rA()�?�4�7#��bٵ|��@J�NT-^���Ш�4"�[bO�Ȣ�Ao]6�bΟkSR^H^�F�������^PFS�$ϝ�u�8xS
P�ɭ�֕��#O���������8x�v����Z,O潍��K/J��4��5�e 0���>�]	��3�����)�=y���'xl=�u�?HKl����$Id2�x[������|�B[deS�n�����W�$nZ�����]\ʝ��k�]�q�vR�z9�
�/�\S�!���n.}�{eSM��%�s<_��E,<�F\���<������@��#�݂2���^b:���֯ CP���(0k��M�]\JJ�'����s��.fC��wk��"{I5��-V"ܥq"��̐�u4�Vċ����9���#��'a}~�&�f/�W����! ���͟��~pl�']F��iS�\	NR�,���� Z����4~�99}�ɿ�)M��ʷ��UV���ŉ�-gT|~i�^��ϩQ���|�W�>������;	/�^�$�p<����W��i�s�����3�\\����V�Oϐ��8��*"o6Ɍ)�J�M�z�\�UsFs���׊}�����.k|P��#��3�����BD��#�w��8Od\s��_������è֗�A,��ɣ�3wX�ZCs�'i1x����_��/Ю��P�9�@bU�Z�.���Y��e�>�̹�O"Tb0'��Ɵ���4�Z�2iݴt6.��~h��(QAZl�^���_}J�����[��=D�p]�jF�;;��eJ�"]����{0��X��R��K,p�]s���I�Ooߜ˷<V�Z0�c�_�$��0>ե�{wO�dX�q�{W)�o�OP�f�t�u?���bv��v�w��T��ꈬ��V��KE��;��S'c*�oHld�$�㇫��"��=|�Q�dI�UOj������ �KD.��;v�?�k��kw���
��F)��s���2~�����M�AUu�����C��/����O��@B_3l�X�4�!�D�^&v*\�0cK�*�5~`�h
�	"�P�EK"�;;M�ײ��U!���f��.�g=PQ
Δ����Q@��I�V>��AA��%��1�7��F���#�j�U�V(��4�(oS�F+�MG�\о��Rϵ�%	�ǮN�@~�r�'TK��f!��X�,O��X-���Q����H�8�I/e�==0W�j��3)�����E���q��5���*Jg��Z+.�K��2O�@	`���g���!��z	��Q�c,�qjj�����n=��7�yoQ֝��J�����%��+��Pk�`Ei[��&�E)x���P�
����D3�ko=�0��zzJz�t�'�ǿ�BXգrmo3�؉�S&��9��H���;�^��9����k���%�/J��k&dB��:g�Mcg�-��8z]T k��,��F�JW���߷m�ۋ2�sE�w)s��	��\��`�Ì�D�:.-$�PtA�cBc�<�~D���� �ڗف����x��oq�K��U/u� o�(�%X�����u�ci#������FdZ�!	^ӵ�ǁ�@aC8즮�n�r	iİ����F�"y��?G\�7l��
AzDRm(�ܣ�T����7x��ʇ��^�I�<��T�y�\ءlT�[n��??}
�o�b&<�צ?w��"2�8��~[��Q�P�2)��7�� �<W�C��]�#���-	��OsAg�`r��uz���jB� y�Pߞ�zy\LE�Я���+��r?>Im�
�xH��f����%a��	��<U�$�@X\4$(�k5�����L�҂m󐱢�U��@�J*^��vi���� N(Q([ˀ���t=a)(��NW�aU�]VSS��I�{>m�D*c�������l�S��*���#�1\�ğ2<���TW��F���R�4�m�@LI�š���t��M�k���'�67�
UM)�����-G����#	���f�l;gT4vѳM�*���ѳ�DUV��*n@/��Ӛ-�ol���7G�����'I1�)���aP#}�\O*I�<%��g>�U�O�{Z�6}�l�K�-�T�1��ί��ȷ59ʐ�"���l�H=0*ɷ}���60Ӥwe�x@��� ���V��B[�h(�2M�sG�� �1���뉝i��"H}��$�*�q��.�"�Ϛ���'�/����@�O�򸡳�TAbm�"��fsscY�{,�H�:���(���9��%�LH����A�6<���N�I4���SK��H-���N�{��HZ�bR+Z����~��3��o���_�9�zX#��L��Hg����#��U��m��7*\Sl{�o�N�f��N��m6����j��Qc�8W!����g���Z�V�2$0�5Q*�#�X!	�0�4 o���K��椩�5"�T�v���SQ�N���S��	z�&0���M��������q�3hX�[��j$ڇt6�ʑՏ,���fѮ����{b��x��7ɡܷ 8��#o�����w��F�ud_~����3Skɟ�H3JS�|uưgh��6Խw�ݥq����>V֞V�5�{8U�޸�!���X-��z��[���
e����T֨Mi�Z���s� ����Zi�'3�2���9^HD����?7Q�q�3Z!<�+�k�tЩ�@KF���BghS���I��[���H~����7.{�������M������>h��]�8�|�9l�J_�����_����O?v3��s1N�T��ҔZ"�C�p�x���]�e�[����i�E��y�#Yч,d���w�-1��O��;A�U��!$9."�,[A����{����>̪-kHd��P�PC�W��c���Q�����%TC��7�k�����j+üiD5���+g��n��^<"�"��ƆDNEq��j���Fߐh/'�T�0�83���u``9�����U�s��ԗ~��wErm,�L*+�%H��#5"vh{v.NR�Y;�rm��1г�����Ɩ3����Yd;mA�ސk��PW�j�*F,��-,*�dRE2�J
���5'����@�3��B�˫�,(oIi����7��m���q�[�e�fفc���_��H��VJLFJ���uv�Wj^�I!b��W�	c�Fd�d�+�LG�$�d�������HHQ����f	���}.���x�L��eB�|��:����*h~��3�������|�w �oe��Is�¦:[_�(*ڷ͢�x|�T2l�T@�px=�*3�{Sb�������pi�r�Y�s%P��=�|��v��ݞRE�Ӏʜ�;����CTD
��pwz��9~uY��]�lQ~x<����X��X�Y�I��V��5��
��3���ab��m2C�Q��2�N��V����Y����	�:��۟C@���Bʚ;�K����g�����EXZ��o���i{�:M���4|���蝡�d�*A1��2���^g���r&X�Iz�%-p�FvE��F�RO�W�Fvk*��z�����&"����U$���o�u���|�Մ<�`k`�<�8��x<�6b�F����W���3��h�'$)����ݾ����A���䐝?-�/��-dH}��U���d�Ks���; �-,��_�Bk%��c�p#��B���{J� ���NX[ک$f 1��s��� �����o-g<�7�Ӄ�֬	#}�i�V���ȢU�2�xшE��ԗ�Γ�)���^�2�ඌ�Ğ)B1采ze%���XK�%Ud�#��a��%���
K��s���5�n[ߊ��j%ꙹ}T��oO�磢��*C��8�_Q�U�(�o�ɔo�r���36~�At,��1��]����%%z4~}��1o*���C��O���5�|�a�	�}�eq4�QJ-��̝d�N�1�����W1�-'�N	��(�瓊�R��K��g:
��k�ܼ���ZO�BSk���ĕu`�Μ���
Gߤ�8��VH�a���Ӷ^�/v[�/Cuu���X��2���� ��bWg���?2lX��T��W\bIk%���7�w ͋z��^���d�6sK{�M���2�z���o�.�f\#��M�z��aQniz �Z�jb��XP�+�ً|U!����b�D�~�&[9vb�8�\����mL���?��~�*pA.�F�U������M�.������b��5�A�1�p���x�b�j��־3��c���Ty�}���*�I^�ʫ++V���i���\F��r����aƐK��z�R����R.��7g��QB_}�		+�ͨ�):�a�f��l�����a˵� 8b���3������+)���q���#�]� S�ҚC����\��ar x����HTR.wqz9�t�ގ_�##t�	#"\Y�7&��,rh^�zN}V�)�ʵ瞛D�WYo��=o�>�!KƧ�4��U �M!���I}��׾W��ܩ,��?�0��̩P�ǫD8$!aX��ޤ��L��Y��i?{��Ѓ��v�*
����O��]�b0�r`����>ߖ֮��+�(���}fz���=EƝZZ�o�_�q��ˮ�g�貁���[d��ȵ�)�b���K139�FYP3�9ZzRmN����"��}�!�tO)=
�If�����t��N��B�� ݹ�0�'�T|����#5��i�n#�i�� ־U��%�X=���2�L:�=�R�g�VZPb��Y�:4xq�n׸p��/S�X=#sU\�x�)F_�./�`?��f$���qw�?)"�Q��R�ǳ�8ڏl�M/�7r�ؾ�9i6�u�5RE<m�M�I��6w���j̚b�![�K&�ිNQ�X�`��*���OKs!a;'�?� �nYW�M�o��QX������x]���r?]�4���{���ch\)�'x]dV����<_�6����:���U혡Yd��<����?y��瞾�m�ƅ�0	��Gޒ�(� n%�G��D��+c�����%Ql %)q�Ғ�)8
fRr�����Q�u�'nR��4�Uf(�����r�[�3���H�S.�H����uJaHu���'��ڃ:�P�ž6pH���T|�!�j�Q��:��"ʬyV�h�ɥOdn��*m�h��~1,����Ry���%C�S�Ԧd��T�������S����a��y�w	�P���8����¹O�8%E�9$oTP�]���<��w��:>���9I�*>GSp�2%4�xh��1��z)�Z�-�Y��MDP�ZCG����px)�S�L442Ut�dl�t�хd+�0�v�Y��H5��_4����_�Xu"`$�M��NF	����H��M�ֱ��:��v\ `*X�'��l�n�+ۋ�����`L�2�m,�pE�O%J@�閻R%#�&��l��W��E.V����5���u̾O�|9Z�H�l8��?�(�������Ǘ����eǋ#�ۧ���/�,�s� nR��j��y����G!�yP���S@NT)��HY�ٴa��30��qW�J
8����>�?�WJ.��ugg�N���.�"���B��5w�[�{k�鞶O��':$-�m����Z��"��>�҄�c؉y���VM�W�y.�`������|���	�\�z$j �:��͇|Vb�d7 �_Ƿ��x-��n_ο�&r�C�)�Ӯ���rr�L�-�b�MS���	���~�v��͗������\��l��k�͓sI"_�W��WF�����R�Ee��L̍�-�; e�&��௴*{qQ�ԫrz£M����˹���򓀋]Et1�Oʩ>}�cz�_�����F����b��5��� Y�yXI9񾤞֠_�P8%���n3���Ͻ��}�|֠`����#G���&Y6�1j�M�8哤��:����6����9��|J�P�c����I����J{�X�,�G.dΥ�	Y�wB��3Y�v/�zs˫MV�V_ғ"�$��5��31�}��9V\�
�t�0�~�פr��Y�v����k�����jP}�7�����4&r��$��A����gjV��Z�|�����*�X��`�����9�z�@E���o��ܠ��1BM�����<���i�����ic��/f)����Ri��]�Z܃�.OZQL�� ����0_)�w Q�̋�~���z-�Uo��R�|�GS��)} �Y\<2�B���\���X%qAtr��u6t�v!�{(X�W�S~�N�v� _F�E�75K���"�zw�M6��Gk p,Ų	�4f��D	��7��֮͜ް,�T�O:�*N�3�r�/��x��zh��U�G5dU�i�K4�H�y��~]�F�D�\�5�"�(��=<���.p)_��M�.k1M��)r`�!20�kRE�ő���K���E&uP�-����vN�`,���fu,�������	Y����4 �hw�Fig�F���:�A����bJ����4��+���?��}|¶�$:<j.�n�0���_;9&�>7řPh��|��P�cGv�S���Q$e���X��{I U+����(�-V�<�WW�����.�������4iz��٫�߫�3�,� )���o������&�@�ޗ�6�u)�zo�\V��Av�V�c��	UjM��CާI��CWN�� 8��&���XR����,]�A��;]t�tS���'�ʪvW�F7��<<q��ǩ�,�4����$����w0�N3�Q6�)hZ}�.iR_��K���rߺ����y���d��P>F	�D6:�ձ�P�Ԕ��f=�mW�.6:Lcl��!K�.A�xTÔ�AB�� ���i����M�����w F�ͩс�VDʌ=Q�9Nt���M��'�R�iY��mRܔ��ߕњ@�D:һ=^,����F젅��4�ӡ���ۢ���*,Y�"�<��z�(��wG��l	���_=�׋��$��:��� j�:p��}�����3p�Ȳ�s?z����H��	�����EH�d!I&���o��z�����D����x�K�ǧ�p��+ ��cN��ʙ&�����S����1Ze"�#�c�M�4�<��.��ɗ6�A��ֶ�#��c�E᜝��]thoeͷ%`Mz�
g��k� ?g�0f�_/&�j����YY^���I�7>#����V&�M�|�oF8�N����An�uW&��͎�N�|��{�
�.�N���]�r��p]���2\��p͙��O@?w�ҍ������2�Qo�Τ�.��8��Ł��dǢ��JW�.��s��>������9�Uep]T_����KN�|W�hz�We�:�}s*ğ�ĕ�wH��s�/��b�Ls ���]����#<W��Uq�k�O�E�
t��V�&�ř9�R�)%���=�F���;D���,�s�O��E�kc����T�^�V���_}�5 ��6V�e6'&#&%���e�r�Q}u���|��f�E�^�U4���d<ZJF�����sn�E���]�_�V��f�࢒�����%�r�z|�P�P��,�����)��}��6c���F\n�k������u�m�;��hy�7� ݙ��.��g��OGTa���z|��|UY�K:�b�e�z�3�X��ݷ�ֿ��6)��Y�؀?x��<�\��V6��6��Ip�T!	:����?U<���Gں�:|h���H\�&)����hTe��y  e�?�J�hB&�;vQR�F�tO0Y�l��~q��[C��77"��t��)��ޕ%A���GqXqP�*c�ة�MX3N��؛�~���$��CnN;%��4s�Q��OI��n���f� ���d"�uI������ˁ����EUO�?���l'�s�ɷ�:xs�e6ڹ�k�+Z��RD
݂h���k(UI�h_x�J����S+�k��zUu�ο�s�Mz�j! �]��~)F�F�pܛo%é5��P�*]6I�����*x\���@�Xs����O���K��E��!w��w�d���K`��!�Fw=��:P]D�ؽJ).�h	³3��!KX���%J��k``���n���@�)d"Kw�p��*cI,��l�h���Eu�5I]O0�;�pL��3���l��f����s��=I�b�%E������C/��������!}��b�-C_=C6�P�g���4���>G�'��=�jr��g!�k�IZ�v.<�ܲA�7Ř~�'	x�x^��A(/�V����a)�h��]�˜�e�%Q�0��V~ؓu���:X�p
� j�U٧�	���t˺8�M��u���W��f:�Q�M��80��k����1�L�c��i����0}�@8��o��at������T�_"�����g-GҷK-S��"�^J�.Z��A9��EK�O̫�e� ;	�ڦj�u<�E`�ҔiC1��`�Vb�Z��\�����O�m�'_�"~��}c����m���#-�y�dy�V�ռq�����;������w�	Cv�$��ū���,����@�څ	�>PX�+��G�e�5�it������?����=�6{���5Q��S9�9���ut0ӓN0��	��n!�;U`_����O�Q$��T�	�,e�\��gĐ�Yߋ������h����.���zGH<���\��������[��
K���I�$���l�-���o�~���b@~Ha��g���W�#e�
����ly�&��,�vj��WZ�I���[�R�C��8�'��W�mY��>%3K�R�\�(f^|�����ڐ��D<�_9�@a]ڪ�	���d�Da�rw�+�u�Or-�P�L�8l�����>%�uk���2�[��1D��L|_:/�}�x���?SDzsP<�9?	d�`�h*�5@;P���%q��\�����.LoB����}{�I���-�e�g� �ۂ�O�:���M�pB��55�Aİ��1�����/�;6�-�Ǧ�V��f��Me鑜�u��q�u��ݘ��F�Zn�?O-�%�e��:�҂�6j�q�N��?�'�#A�]P�^K��X!��8�zS�S\|ܑ2�0��#�b`i�Љ5�/�I�Ċ�G:�}σfNl��?"
�vdo�J-E� �f���)�VT�~wT���S��w-(���m6��%"?�����ʱ�2�C��{�KK>�|.�eO��z�l�(29�6|0� T�8��R	�%�3����O��Zzi:�1�SYrܳ�r�0(M�%1�\��Iİ�]�(�((�~oL���"��Up��"�(mŝ����w�?��~5����0!�ݬ�*#m�jٙ>�r����EN�E���9��g`�J�vq�]:x��q�i��V���ݫsKl�>����NS+�Jv��3�?6Ry��ļ���Pl�K^���3ʨ�q��6-󔑂�e'�^���1UUHGh����� �!��9L�5��+�-�C����ꊃ���X�P�ww�8���R�])����wwwww�A���?q�m.r�';k�$B�t1�Ό��d�s��a�����_�;z� ����C8'eG+p�K����;X���M",��n.�7���l�Ȑ��1�Uȴ;�+�Sg�~������xt]4�U�Z�W�z��  +H>�R�5u(�HPu��*�Z��F��m�k*#�a8U��:�u�2`��K�L��NKco[�G�?\�}���zm�E���Ʀ�i����%1�N}ɔ��鉧����g�^�Ap2��2*��F�Ьfw����Z�����[����1�Rkp�w��W�^��U�\=��,������j~���l�L��{��숴�eH�N����������H�X�,����^B��P���Sws�S>E�@T�S��(��6���r�䩻��8?���ְC޵���'d�=�����eF ������q4:%6���eZ��p�*��%ȳ�I���e�f�oKe0$��n%*`b3��<MO�h/%��+g�cW���%���_
"������ƼK��m��l6��:�� S�nQ��3��^�T�<�Ź�<� �y�Ӌ�9!�|un�X����r����/���`�4�������v���va=h!S���n��f��0���9+}p�F�U�?-I黪Ɠ�U�EM��p�#�wӵ��l���xDi���rG��b0��;Q���Y�8tA�����Qp���v��l�p�o�v��ǰa��qt���z��U�/?�Nc���� �dO��ed�awҾ�߮���ԟ[%��_`}�a�SC���k����]�*"��T�qß�Aj._)�[��$��6G�L,��1�M�����z�K0E
�������Waf@|�]�_�h�}o]/LK:PO!�O
��ڙ�4�x(���7x��d�8i���u@=��vng�Y>���f\�{��}��(��BFe�P�����\�깦0�cJ#G�C�����͙+M�֧��J	u�Jajc��r���3�n����#W5�����~�)�=��<�m��o��1��J��\��}x\��=&YZ�`ˤoƳ�׌����V'��F�.�I�W[�<���+Qۈ'��KB �u ��K��z]xT.��O��M�HQ9��򰄺���{�_l���A�oz�m<9Z��.'�֝�R#"v�*�m�XS2x �b,�x0o���$�h��ȅis@!���J�Ή�

��U+�V>����ӭ��	s�_��-�+mg���EUQvt\Ը��k�R�h����
��\J �Oo�Şv�B�n��!�����=Av��C`d�@�[����ͱ�iȤΩ^M�P�����|y�ٱ�ms����u���{e�5G�Y)��
3H^�n��Qs��N&K �R��Z���~��fT����a���}T5�7QK&�����Z&�{=:�ǲ4�����B���6	'���h���@��aS'���Y����{��'�#{,���Mq�0�y�W�;Ƶhh�_Z�ޡ�A�\��oV3h�7&@�sjm�EŶ�f�K?zgM��!���v��S�/�8��㖊����3���D�U�֙���n�U�Bm4�c�-g"�N	��������in����h�ir[#F�h� �d3/PDg�
M�4�·y|f�kTV(抝�%�����]t�RA� ��F��%M�-�&�V��ZN�[�ұ�]�_�G�.$�JF�M��f.�q^����8�ɶ%��@@�qʾ��r���0��߲�����פq]����s�4ibc>ݜ�>Q+ջ�i�_8>����C�w��.����ȼzk�q2;���Z�Ɣ.��=���� �!�9�����
5UT�&��*�T}������(�八��KA��N�_jwB@ްEk��(wL=�Ѿ�+r����&�|�UW�Yq����U+���J��~8S�������B$�/-�<q��"6J�G�����I怟�Ҟ$�y1�0iʘr���_� �֥�$�{,�F�<ʋznUk1�����ش7��ߵʇ��7V�W&�1ӊ�]�,�?T@N�����տ�~�: ��Op��Uۼ����\��@��2R\���D�0�}�XBk��~�.�:�%�7������16���3$�9%�?y���D��!�xj_��X��%a!{m��VϚ�Ԭ�h���� ��w�/xg$�m�4�V�9��/��Wof�b��Ml&Gj5����G�U#��8_�hy���c���z��\ib���h�e���(tn��^�pP;�;w���bДS�uE�[��7����.����)-���'���L�o�|��2������u��=��[@�!���ɚƕ��ڦLu����J�(ר샂f�G� ��3����̛��f{�\��棩����
���\�Sm{�����:���><������W�I�.�NӶG{V[��P�ϋX�%BfU2>M+�L"��R�F}~r�����X'���P9E�����eV�i��!��=��2���L������/͙T����-��Ļ��x�4��E_���&)Bl.^Q��{�幔�����
�o�ރҕ��Z�˳/����,�;���5L°�3�7�֕v�vM�A��ѳW����	����@A,K���hgi��VN�d�O�h郚��",�p��OUxx��u5�&��FvU�+</܄3���Pڇ5m��+�Y�%��K>�r"�=�l�+q4�`���7�^+|Im�/��YkFi�bT�^�˶1�Նq/;4Q�T~���0��%���+7���W�Ht��ښ�ģ5xEyeZ���(M�p�xgJ���j��|Xl��B���;�e���)�Ƅ��-��w3A&x>�d{���W�s�;�UÝ�@;ܤMjALpb~�_l�?Z�=�%e�¡�i�̃!2�
��Ey�]�����r����E�`��E�>ˁڢ|=b�d$���쫲��I#Ӳ���
��Q,$�ck��57���zFb��˧&]�A}뵾���+:�h}�a[>�Ó�6A#���I�hȈ9B��3�������9'����|�{��cO��7�kԒ�����C���/Ƥ�ko5����V�\��w����s
ڔ�b(d������b�R����@�%�&Ke^_M�{X�0aUd���_�TAI� 7G�Nڅ�F�a]!���ђ.��e�+��俹�t���NɅ݊�1`�d�~��h�U��dS�z��3�R�����) 7��G'6f������v/����	&#:)��	x{m]},l��)��|�i�����Z�R��/��H}RWlQ���k�?��X
�l���Y�jl���x���c� �!�z�ln�sz����L���d2�z�u���-��S2���[��XE�֍�kE��l��U�zY��"X��g_`�y�K9؝��}'!I$� �U;�r�z8����VieFX�F݆�a��uh%���__�� l�IsaQy�<*���ʫAHR
b���(nz7�Wl���z��h9E�8�(h��?ƻ��VR�&�nN��)��Y��Ү�B
'{��&> =��#k.�f��Oe��8�F��n�!�]�ߺF���]�j��GY�f�0�V��M����Qbc����X3��)�>x6l�m/����v�O���ey	����B�<�1-B5^n[���de�Fޙ�1+���琉���v弿:!N����j�u�LG��ʥ
@��͉����R7�u�b�2"a�Y��d���j�m���)cQ���W|�������}��~��hƘ��f�l�D��V�,����&\���H���^b[�ٖg�@�/Z��q㪓�s]�����u�i��g|���#�g���N�����v���w)�i1��Ys�zŚ���:�H����2ϊ_��=�g+iPV�S�T�A����T�D�{�U�KtS��Q�c�#^Q�j�tLN�`�}����"4m�a�QCrI��o|��@{z�WvE˨��s���DW���}�Ug��7�[?��$����>sS9��F}�/�ٚɆ*5\�P�����σ �`�)N��ҙ+�t���A�B<��^T�7��'K�lm� cl��;�&Ի㋑ɉ]��H"�r<��R�:U4q���K*qS��r�gk���a|�&�.U�������ù䆱)G�[-D���A�ټ��O��d|�"�߅�dM�Z/y��N�_Ӫ��	�*��%=���i�S���}"�@���**�e.�PyZ�c����+U����wh��Qk�)���UϦ���jXkt�2KP�Y�3�����^
��K��߾AB	Ir�y��,<�z9�Y�<=�/�W�v<�-`8[�+�ü U/����˧rש�1�y�|̾:/:,%k�����ʝ_b*�Z��T�$ҟ9s�N�ܴnt���(�hR:$G(W.��ԡ�Ӡ��`���<�S���?��]t���	e���8�F R Y?�R�e�{�
�����|CΊ@I�b�V���y���,K�8�Qjo���l@\#qy_);�9:c�O�"�4��H}U���D�?���R������m�44W�[�&�׿1�ȿ�:Y�}���sm���\>�Tg�=[?��z��xȠ}���3.jק�٭�	&�IX뙚�ٮRBr*�)&a�����k�d�D5iX��^I��ϝ�P���


�*��@%�-�]:���6=O÷'26}:k�/��<���"G$����d�0R��!۶vǊ��-��_�?,ܽ1��`g�<ܷ�K|C�J��h-��>�� pkX���bi ?��|%�V�K��<6>/�\L���j�%��N𖗝�������BW~��U�E���drkg�W��O��a��MA��Z�ߧ�=���5��Fy�-��'x�6%�:�r�Yi��Y� �����2fmm�|G�@��;ϲ"L��&%�Kahth��hCU�����X�H��$��vG>͟�k�d���|'Y$��<�:�k���ȩп�і���h�HJp�ڶ.Gi��~��UlU�GwL�p���/]`���L���Hb�6mˊXS�}���HVܸ��{�ݘ��H�DhΪ�[�uMN��ꑛ����.���?� Y�gF���T��QQ�a�� `�m����\�v�Q� 
��~&r�]�~o�/w�:�0�Zg��d�	�%wKˇD�	�4vCz�����LC�����F�J�W��tl���(b��P
���F�"�3�"���U�1 _��8����<Qy�9��:�*
�T]<�,0j�,n�`�-L�`{���*vB�F�c&���c��g������OD�K�)8������;�SG�:(��(P�V��t	����z\ڏ�I6���3�J3N4-�b���f��k�i�sf��3��0�@���f}�z/t�r�$:d��Ei#JYs��:��
�H���|P��ƸX��}�Lə��H��͘.ܴ�Y��]m�e�+�p	��z��C�F�x�V��OWi"ø]m5�=4Cc���Y̵�C"����iG��Doq�L�_����;�>����^��;��~��N��qǻ ���c�`8���3���+��@�x"�]���a	� 8	8{9�Hf�g�� .Y��P��Q����5�j^�V�G�	�!
|D��A�PG�9���?�1�S���~�8��r��%��t�a�����IK� I�]oO'�Vץf���R���#N��K���oa�ĥz�@��f�9f���{c���(��/+����2��v�ӆ�D#���y[��#�$�0'T>���i�\Xsm�f�=Y'��dz��2����7H�f�V�>�s�*��(�GD������XOZ����ܘ���٩\���#�tn��xP76��C��ׄF~P~��i��Ȫ)L��D��?ϊ���;������9��5~͇��r�Ɗ�t��Đ�z��mx�?{�=y3�{�-�i�����6�$�!������;�ß���n�y� �?!�����楼  ����d��U� fq����Xx�<�X$Ln 9,��(�����pŗ׉�'���LǈԮ``�d�=��J��ΞZ"ne�h���,���z�%)b��X���>�߬�]J ��\0ko�q���jQ�z�^ϭg�ʤ�x
��͢>}fn'��v�8���ke��.��Z�Vꨞ±p��c��.��d����Чx�u���LZ2��֡Ow/�ԑ;�_�����!���x�E�r��qs�mb#<����[��z�{x߃���}�dC;�OH�1�T�e�P�U����Ji]��=����<8�P�{���a*�S��믹w5��|6��B����c�ڋ������Y�P��Cۇ�y}d����K�*��g
���=kK�� !�-v���0yK�}׋18m8��m���G���,�c�i����-��Uh�5��%���N��~��[ƥי��&b`(dO���C@v��!q�L{s6�i;0�G0u�+�F�!j!�\�./�6�
*�"���)��MtǅIi��+8,&�,fR	Ű�q��^�c4�X���J=���"����M���G��شN^�$�Kii�t1&��"�}qe~��$Pk\AT>��"����2<QY�І���`�F&����92[��u�:x�����QU`5k�@������}���m@ΰP��u���Hd�
4�fr�Tyu�)/�����%�Qn��B3!�	��H���7�U^�aߋݱ���*��3`n�// h�OLiT'��-')M���v�̯�?�V4������oS�/��vC�y��c�}��>T)9�.�l?퇩�g6Eٕ�z)�Toʙ����ʨ�qLauDM������"�^�ܟ���.�l�c���r����A���D�a���
��cd�{�M��{~/����H��g���I�S��4�C�'x}��=�T$���5���E�u�_@�Ӧ�|rRB� �rq������VCL$��`�Y>��59x�	B^D�P��(�T����M����SRI�1���0���c8��{_]�Q���Ų0]��`�����N�i��Rϙw�+��]w2՘/>��㼎0�0?�s@�dq{g��?���bxΰ���c��ق���Ae#8y� 8
�A�IM���j2���]�mo��uW�Ś��D���Q�]�����>�1-v�'	���r�N�<��ؖ��T���'kR��&YP�O�J�'H�V���,o̷�52$ݴ�0��Y� �s��)͖�>/V~TdFs9�H�&s���2�wL��b�y��N��1�I�J���1���V�,� �II�G} ���ܧ���~RJA>� ;��	%&m�\�s����-��Km��m6�"q��f����!3y)����(;Mq�o�<�f�!
�|㇌��e�r��:H��	�? b�QS�P���Z�ąY�#�ͳs����&*�*��	)���a*K:1�)��)�	��x&X�5k��Ld��<��n��QULK�l8*�^,��%�$�#���/]L,�����4\j6"=��+�x�H"5��⹺ZOR���tn䨗�m�=\��е.�k��{ �Ei�>��  �_~�ju�_W&��n�N�C�]2��x��9�$����K0�gB�v4A�B >�r�_;��wD�m-�|�/�2��ÓR�ã�e߹��^#�մ��>W���	�0s�/��g�U��#3,��o�����]SY��m�q9�������l��0g�kf��Ǳ�S�]����[_�X`��`e�;�:&��c'#U���_���w2��,�+Y�տ����)�^8���G�i���^�^��-?��Pk9gC��@u:�.+h����u ��kT�K_B�R��S8-~h��y����R��}'���׻5i���~��޻�Jf�ꨡ��2��(~x�7���=�8���a-�$Z���@�/e-�҄&�H�%����}U{�8�0t���v�3p�ε*��p�e��`��P���TxK�Ъ8P�݀���T���J][�%�:w��j7����˔��I7>�ݷ$������/��T�����\\
��R^��<牾9zpJ2̎V2h�*2f!*����j�:r�lǳv8~��i(N�_�D�*f���c�)4\o
�e3.��u�܇x�-�ߢE\0��D5��DN۬�%��YiG�S���:�}S�Ìu�w�lk�X����RV�G�iT���t��]e�Lz|;��|����WV�**-�E��CJC��%,Y��� dߢ�F�Fe��֮�D�z�#�YY����対���4_�vk԰��I��8�4�c]��������=��	�-���p�Dmu[�(�Mjb	V���rI,g��?�G�#��A0��������w7�ؓf��&x�g��+�$�4����R�Q]zb1�TW�]��8T��r� }�-�����w҂�}����(��uv]�3}Gr��53W]��Cz���(�)�$K	C�U�Ԟ��ND>�����h}��Z��V[��载/����	)o��|_*.NB�ըz7��%V���n�'���S���/�]]*�'GHmH�
#"�nl!�[ȶ�Du�U]��5��~ j��=��A�,�/�И����E���%ړSrnx��Ƌո����?��"l�4�"��Gn���������ݰ���S"�R�l���0J��:��o���;�8wxɉ����.�R�h��)%��0��W�␳��l,�r��F��"��Df)�f	��s�h|��#�%�f|��lnطg�2a~�EE� ��b(��b�k|��ZpԆ�˭�u&E�c=�����~dࣩ%�����/s��ȷ[��E��cߚSC�O���P��Z���g$b!��e�����h�QGQ�;f���s��9&|Z������jR
���z��V�`����L7�R�WUzI�=8ϡw�{r,�w�!�h��J�|A'U���k�Ҙ���^���a�6����L�b�[�A���G>�q��si?Q�Ó�_��nE�Z��6�t��60S	ۛ�S�"]��|�y~�c�tcbH����KD��&#\�d$ٚ��K&�Î.x�*(<�}Z)��l3_��K�
�{�kȋZ)�m�{˕⪐Q�*�"�1�7J��+�J�va� �Gϸ95��71;s�xN��+�Gd��3u'wO�ݶ\�}PD5�����Vǰwº�nV�DAQJ��*��GR"l\��5X@o�Q���*��y?������ ;�����Hr�����Y ��M7���to��`=��)�%�+JM
��5�`��Bf�R_�����cl+E���tU�S����)^s!�D���/�V��<�x�>��Ŋ�w5��^P����QQ�����ur��f�����zԹLB0(��hI��`���Z�˸u/ �I��
�����7�&���9V�S�\QsH�{:|@ۼ�T�|_��3��/���8H+�WM��"x����['�/���!�����R�eЅsh�#�)�Ιl�,]}����km\@ �I;��8����}b�Xn1�0����B���Ӎ�>�fn��Dth"�.���Q��o����`e޾��ʚ]t�c�K��eg��y��E*%�:�-]kZ�۾u��sF?���$��q�b���Y1 H��U�R�ZR�P��> |��ѷ�P�em��2.���@j57������e9��u��J��M!u%Y��~�o�^i6lZM:[-d��B,@c�j�v�U9�-��_��3f5�T}�R�B����Gwk? Wq���;?LDv�4;6�I�u2T��A���5=��Da��݂�V��.DN3�����}0�[ ��V�1�� o��m�v�K�P��Z6����2�"H��w���#��� ���|ܘ4އ"T~+��2<��o����x������:O֠�~�tC���Mdi�^.��3�����	�IMNNW�Ĭ��9�Yuh�,�y8�8}>f��7�4����'p/�b�[�a;JLH��6�~���Ɋ_���)#�� �h)����X��	�u�Z�6�L������7.��^�)�/6��neFO�PǾ�����t��X&&v��QGҒ�p%�|���e4M$��ThEK�Nje{tWk@�pb��P��=�JƲ��.2����b+�W�S�()��`a����o�����EC�H����V�X�w���vrM�L��e��^f�&�RA�-�Xm�_�1-��ˑJc�=NA�{Q"�q%	�2�e� M��%�D~�ۅtXA�B�h|���R�q�[s�>�&�hӢU�O4��o�S��~ʤ[�x��������2��J�Q�?-Ya�D�,����w�JK={�V`/�����?<�M�u��� ƃ������W�P�DX�2%Ezq��2��-����} }����O����e���|ƌ�֪�Q-��/���ǹ`-x���!+F^ZEm5/�1����^@���6s����+'�=~�I�4o}{oU���(=۹滊�rߊ�2b�`=՟RӚ0Of����0�1�9�L���m��ͷ0(�SCk�!�tVױ*�����6x�cB8����.|�oDꦦ���N����H׭�zy$��+���w%��F���۽���x�<5���[����[�2��	�5q��Jȴ]��Ь����%3����,�3-���![�2�l4"RF�-I}>yG����"�V&��X�[�c�m��<��QB�i�-Zgs,�]E�<ࢰv�į�V��_bc�~:1Mc ^���ţ�gGs�/���2'�<UPsLq'���@�\\O_hў#,�TY��CV�۸`_���]2�� E{��x����J$(��ɫ1lM.3���B�g�y��0C�{��ޙ�c83�f7���Ҳ�qX�n3`���^o]��t����МnAV�[[�MYCJ�^Q)�y�@�ֶ��#'y-�n�'V�O/�� ���E��S��v�J�2�a��7����n�G���R'ν�/,y_յ^��,6+˼3�Q)͗�����F�B/���d��5�4�|	��Dp�j���C�����@�P�%z1X��_�i�N�0�*��TJ���82�Cn�CI!"��������kD ����7���.�M_P���E��u���	����o�δk�4,K��UC��b�*Ӣ��
�x{^��|����d��̤o9�����׹�k�e�m�C˧³��̣@�=B���Jb��奖�?�*�GбɢZ��|�j��Y��	t��c7�+>�E�HSU˔���z�k�`��k��Rsj��3�Z����<�������
u<��gK*����|~A]#t� <��`���:���\>��d �c�����B����|!��D9{����k3~��B��;B�J#�0r�3�����j���܋�w�����>J���u�"D�"�D�����h�w���(Ԟ�D�%����H�!�j��p�B.>c����6�s��Ka��(�"�|��s���u��(�=��*��w�5t�4tCb��+P\�y��`E���#{:�v4I,�Y ����+[�j�[�[�bօ^H ��E��X�45'+����G�����	,��~����My����ve����[����Eժs�7�n�J����d��=��N*�pc�g�+�����~/l��H4HSBd���<3'/�%r�<\�:9�[�)�C���S-�Y�ʡP���o�`�;�V-���6?o�rG��r��G��7�:a�{߁�(��PY����ܡ�UWz~��%ܕM٦%ۅZ*��!�i�!�d�ɚ4 b��4��W,�"ZV`�Z�!�(����VO��j�,9tS|��z����N�C�2{�̖'X �t��+�P<�,��W�ݛ���Lii4)? f�e�ڍ�o�������Ay_]|D　;t�]i!Y��F~1zaY��V�=e
U_��,N	;����q���q�X�<t�e���f��ϛ�6�^?�6r_$�'sM��.�����`��n\naA�ӑ+/�����-~)�۰{��vQee0��dW���6�+����`���cك�e:�Ű�â(0��Iu΃��g�]��NRV)R=XƳ�4�wW�<lp�diF�}�a�D�CĆ�:�.��F �A�`J+��&��M/� ����9o���zm����D��Ɇ���F~�W�UXѐ8Y���P���Л����W$��I��cǫoa}�(�|�������o���\d�O�(��~;UR��r�e��kN�1�.��� �"$��!L�u��+�L�P9��P���xV}�W������`��T�̝fV�S�V��?���)������?i/���N�@��µv���OB�e`�z�q�@��jt��e�ep �`~�̱��̮Tr�]�kT�fXT��4zb[����Y���c���#=�8=���hȋ�4�	��#�㦄�sx-���oP4�3���>7U��=
��S��'6T�;*|�{���Ef�D�(�9C��Rت,:B�ŷz��)����8>k+Z?����ja98����tpv Ith�3<�K0�k��宩�B��z�['�&|��(�C6:�/�,>lr�Zѡ[�����q`�]��}5�U��ű�T�'�oN�ଳ��d��v]����$71��[����$Ջw��^����%���ǚ׭��R�_J�� �<]�����hg�@�����^�7�Ι|���t?�:�2`$�T�B@𹍍��͛�(.���؆�K��$7��")���Ά����������םo�-�|����(1%����YBOGG/f��������X���s��)�K�L�K���+�>���@���uM#R�#?��j"���{4֧�&Vi;oؚ�����\�̍�L[D��2|z��P� 2�gcB������9�����Ғnũl ����t�w�	6�����Z7.ɓu�W�O7��.�6�5mM?�؟j֤~�ë;I�����W|�(���ނ� �#z�a�Qy�n���W�OM����� ��y����H�Ue
�8��eE��O/<�M��L%�FF�u? ���zgI��ЙT�'���監H���X����.<N��DZ���ySא���ܪ��#�9��jb��G6�LU�x�OG>#(8yM����;t�D��I2> �g��D*(}���s��YZ<f��Ϸ*Y��;�v6S"�8��]Ǻ�ԯ<� ���ɒ�k�	��b%[K8y��9�ồ!9G������ο$K`>s~�=�Y|��q�QfQ�],��O����ߙ,�,������5��y��I�Ų6��a��Z��'}~E�Y��Er��Դ���BɭbF}bg��SL�v�7	[���\hC��T�O��}�|gkw�� �7�u>����J(2@���~�^��X�Rgt]x��ٕ�MHJ"�z����r��V𓄪�K���t�P�̧5��K��%���������<v} ��Iy��K�ԟ�w�%{gP~�Shm����)���.���{k/�O+�� �P��k?��yo������f���q�x���{����W!z-^ٞ��L)�k8#^D���Fh��p���R9j.���}�R������Q��!EZ��L�-$�z�}@1z͆��	WG�D�������|�i.�sڳ��|��½��6�'�>F"/�PIH�ڦ��-���.q
�	�����dUk�{RC7�Rn��+A"���M3�=E����_s��/���2+�P�ܴX���vM��(��V�A��jDX������K܇��r�J�*�=�*�_��h�bS�����?��ƪbMjs��H%G1z��m��EJ�+��@��i��n��
�G�	�
�h�s14.��J�� ��9z7��E7b?�S�fn��wj+H�e<���T��Z-6x���!�XMG��H��I`^P�
#�I����U@��VN�]�B�9�'U�8��x��s�$��Q�o|R.�U�D��;��9��O�ЯU������(`�@̋��&�b�S01��E�N�{�5!�&�k*��1AGw��r�^R�]��z��(b����tdܢ2����}������'�� �X0dŲ_�X�;Z�Ѕ4�ז,jG&�
�U5#hI��-CV߫��4+"�1�+E����CoO�t+�� �y��h�t\��S1tCrX�����9�z��!5�����%rTEx���^D�n����*T�����S�.���*�;-����@�U�ԤtLxV^���4I�I�$c�2͓ۛ��Q!��G�=9�=�hI�]����4�����ѯ�
)��Q�xW��B\���^)j�K�tè���6��f.�~:Fu:$¯ˁ�f��N�o��L�i��j8�IOC��E3�fd5U�jDƕTi��������[��H[�6�j"Q`U��hu�,�e t� �3��W�����>��A�k���k�\�G�s���Ҟ��OE�(-��>hTa��q8�����)̸��Y�?�<��d���˰DI-=¯�2�0�#�׾^�ӹ����w�UN�8��lOo�I@&���5�j�� x���I��`�.���D�6Ad�7|����M��1���M,���Ҕ�C?U$e��^��\��� %pr��JN��ަ�ӛ���~ J��'s�U`�󖰥�]����h��1�ߌ1��Q0_�ԕE��cZӸ[�Y���w+�1����]�c]}6}�ʠ�b,�~�Z���r F���S�K������W��|K��ԃY����#gz�h"��_��}|���ȧ�'a�<���4���|��d%}&oF��z)��9�=4�X9��]�Xv�6��x�$�����VB��~E�������� R�Ē�@jȐu���j�Q���|`kݫ�������|z��?l�_ms�gfg�#rݜ�R!� �uqx��Z�%�6�y�\V/�{9�?�5˱�Y.�*[J��=(8��d���V$�p{ a�תyO�`
B�hIi90���,B��	ك*�3���c��m���͢��p��o׮��X�Ѐ�<阵e�i�	���#�T�$��	2	ء��n�U����6zN6�����A�aH�&��R�:�ִ��iޗ�/Z��w�2���ٿ�v�%7��7	�Q��qyy�%��������"�ʲ��&��~�,u=`���=8�E_�ЀcB��*��Ҧ�|i����E=���'Z<ӫ<����e�4~NGU��"+hʰ����gi�-��(�j?�&�'�qĕ�,,��c;��| ԫ$��dA�������rA���Ϡ�����f}�>|6F�nE~�
h=rrН�؍ʄ������%��m�
mp4	c�!c�p�Q��K,�>�uC�Pg��l1�v��*���j\]]�=�E�F���8����� 1j�"��d�Ӗ-􄻳|S<�,�W��d��+=���	��wT>��?M��/���Q�|$���Ѭү���� ��ϋ�jck�0�*;������0��>���P��%s;*�`0;ƅO+���|�����Ԩ�ł����Ĝ�$��?�~����d�`�(�����"���k���妸S�&e�
.�h<;�����1Lp���0hت���\(6d���nL�*���l��+/�����a	�2;,V�%�`B��X����FJ*��������k�/;T�N�Ew�G����t�{�g-r�k�Gk4�E����4�z�I���T�]N��ލ��I3�ⴙw��O��^�PGo�r�����#�H5��V�n���$����6c)u��h2������2
��`��@���o[��1��>G�er6H�C�BgX͗~��u~����0���e��o��@ژ�y�p�憇��,I&ɼ׈LM�W�y|_L�u��֮|8��7��z�r��������v��pCm�B�Y�	׷|V"Z*K���\Hb�RD�d�W�RI-�YBK���M�:/�چ�����M>�]x�ݤ�e�S�hd隶������yV�^l-�����9��=V�>�,��5t�����$ix�.�/�F�v3�?dEi��e:�#u�'O�m�̠�tY���鸝����B���j�?����ꦊ̴<�6	�4����44 #��Ϣy�CȚi[rj9F��Y|C@N,Y=<m��]�B�t��a�+��նw���Zd��R�ݥ,Nqw(�eY\������P�ŭ�����]��w���|�Lf2��K�N.T��wN�}#�fGi����#�c ��Q&��{M!�����G���c�|v&���|V���Y9�`�C%���T�SbWr
��qf�/�Rׁ�D1��כ�Fc^�W�=P���R��$*��z9�Ah5�]Od��<�����ȶ�7Ck���seK�F�۱M@g�<M�ȩ(k�ܰ$�4>T�������Мp���~�-�ک��l�V����ԡ|o�U�L��A����Y�ހ�\�B!5��⳾^�n��H�����@�%��I���2|2t1���7�Gb��v��a��"T+6�~˶�ˎ�5����;�v�������m]�kZ��Gꏹ�йE*�����q��ϊ�î(��HƆ)���D:�X���\߱���8���tԕ�	�'����&�)��	�ۂ�ԑx�l}���.&��,��tАԎ_2��om����>��"��O3B��V�52�fMY?�K@�>�7�Τtލ.�������:���0�J�Nl�&n.	�fhEo��_�N�=��}������������{Cl�V��Ռs�@����h"��~h(6����M�g�y#mR�g�k츬ǔd��G�K�͋V�w۴-�mJDZ�����vyA'���O��m3�V�[��I��j��r�D�mWG�����?7�#��wO��DD��*�a#���SK�X��kF���ψ4�NQ�iCB�+��ܚ�ճ��BlLİ�p���+������!�3��6��>T�C�U,�߿��NI�O5B_r/v�pזI$���I)�;ޠ�de��q~P��F�ｻ�=�j����ꔩ�T�`��_�����3~_tn+-�q�`s��s��RRRț���;������5��j֚(�vq�oxQ���]�Ggn�\���mmN�C�ֶMJ�{�����<P�W�W��%K�_xxڳ�_M4�@x[�������\#S*+����^y�j��.�Z^����9���ɈA� �=iȇOyȥ����x�4Iݾ����B�����y�s���x=o�5p ��#�f�2���u^�n䒖?�� ���JV��{j�(�bP�`�.�8s�V'P b�9�8k��6 q�ha�&�uGk�^���BZ�6�DR�B���4�v����'�݉�Cz������:"�=Rc��ɋCI���]��$�I�&L�0�������e[��5{��_y��q�h&�^�uC����̔�g��<4�(�|%��^�j�rij��涘I��_q���E�U� In�� �.������Ѕ\�BFY*�&��ƞ#Ka�ũc�Vǁ�X�,��/���k�O���2��XX6֯�- ��hԢ}i����Z8T#���XG�箤�g�R�	W� �X NV!���8?��4�p{�P3[�d��t�-�X�j��<�T�<J��i��@�X�E�>к3E�OP��jp]}[�mn���Ag�;�G���ٕ<����x�9DB�C�J~�c#j�R�v������T8s�xq�̺q�31���O������E�3o������X�x'�F�hɻ�-(�˿XөĖJ�����ۜ�(�`�V1Ub���TL*��<���s�IfA>N�8:��s�g�>����кus�ۥ���%S�Z�<Z�v�'G�v�z9G�L(�����Ǖӷ�zʺ�<R��ץ��_?�W� հw���I��Գ�P�}"�cym|���A=#Y�_}�8�veş��Yo�t1��@�w�ѯo�����1�,���>�?E��QE����!���
���9�/��C����G7�m��_��>��������Ơ�4-z�A~L�~�X�'�Y��	R��M"�6���}SS����՛����`Q���0]�y�g>�S�O*�f&����h�)Ԗ�c��,c+wd�����o��b볗��"��%2`���L�>�n3Lmm�+�5Ҽ�̚[�e6��� �yA���k�\�w�^7�.I[�+-�3&�Q�Ej�0mz{��a��b	�sEiD�
S��\��`Lq�F�Vg�͕�rtA)VSCFM�h6�q؋�X��xծk�.�9n
[m�&����B�8������O`���8⴪�� 6A+�+]���)~bVI�T�Me��>S�r�T�6y.<|zP���+�N���a��a��������Q�O�g�v
��=����W�!�aEJT�3υ�MzXm��SV�Y��_x
�)��[RJ}x���9�����oe��@��y�OWI�^��0��,}�h*E*9�V���61��J#�L�'iV��;�F���c������H���S���(����Ҥ�cƯ����B%ة�*[p)i�9�-��ͺ�q�&A��s��c }�-y�Ck�C�VoX�1�&&�ASz��qh��D';�0]�}XdY�N�g�:{!�T�ނH>~�g�*O�I�lX����.��3����!�W@e�a����])f��}���,H\�&���7�I@��O[����^�q~�\�����Mo5=MW�}�jq��%�?,���	 {�-����}ý���E,@�01����}�ޓ�������M�l�eg �Q��Q��Ƈ`�|%_�
�x)������)y�ɐ��T�u1�Y��ۧ�,�a ��C�ؒ6�D��]ߌ���7���:���Ȉ+F'���5�T��%�)�*�J�S/�'\�w`-������e�D�r��U�cu�rMwb&���\�^q`�T$��G:o��2^�������w�}R�h{S��P�����ĩ�0�
"�5*3'F@N��o�Y�w=�ۘ��) p���T��xG�+,�yJ�F=�H��OO/�Ŧ��c����Q8F#���+Ua/IA4�zHM�������"����+ �t~N�2>���*00�p�������+��"��Kя��+^��H�?��<�B>�Z(qB���d��TKqX�����_�(�C�ae��B:4@H��gƝ��B^ދ����
q/lgj�F�tX���-����Uc�x���[@ݭ�K����	�GO����K`����o���Y[�D���@<ɤ����f$+<��˻�Q��u�E��L�=��J�k�h�r�(iZ|B���W ��!�x��gf(ux�'�4�͗}�y�fM-NĂt�� 5��"�X��'�[�c��,����%ņn��Rϼ����Z^�|��o�~s2+���FG����I�ʣ�$mҜݵp"�b3�:r�닂>��
WC��P<M���x����V$�u�:�ퟱ^�mK���=]#���6�a_�4���??��N/�l��)�'٤��rIP ���.3��j���-0�'pyjy�Z��=(��C}Fc��tصfC�R���j�y�[B�p�l�S?�̬���
`�a��k/|K�mtKD��H�!LJܝ|0K6�j��9s��{i�.Ӕ�K�Dٗ4s�䮼n4�h?g�p�����<dfX]s>χ�Rv��I/�+�i%!h���a�OFG3q5tf��Ww�?�1lPQQu94���iq����^����CpmU�E��PF_�R��''XE)&��5p$*)C�%���k��H�O�j[�%H=���^u����
H8���~�ի��
P2wy?�dñ�pJ�u�@�%����;��`1�疧2i�I[ �8 x��<J�;Ƭ��*����>���A�ѓ`.b<u|�8f��q���Փǟ���Җ���Q02�_a��t顉Kt��R������ϛ��F��KɁ�?㖕�H�����M���H�g����7��ĸO. �
W,%+^��F��S)�h��ɬ ���X�\��6�8��Wf���"m�/<��L�s��P4J� N��߅D^���P��^�)�����N��\H������QI��d���s�����s|E��l����Ν��8]���?�&O�����{�?���D$��h���8Y����1���Hb�2������n��>al&G|	���z����Q!ְ3��is�����
�m7�E�І�ɜ��F7nk�'�Vɮ3�y�W��ru���	��l�� P'C�����t�}�$+�%n �bf��%����:��ɶ[u�Ż�ڣ�H�A���WO�"�c�X�O�6ͥ5	T�:
\����*>S.�ښ�z<��������kk�kR�VG��Z�ؚ�9�I���=�F�.� ^�����8gp7�\�؆�Q�����n�8ǚ�7�4���˗��R�q��"�uXa1)`,�E�Y�!�"����+@�����>YV#ގ:��'�<��R}u/͢J{I#�$�tG�b}�hrzat�(��(�h���ZH~	��c/�?��v��U�^<0�h�	�!���3Jl�2ŗ�Q��p*�a{��Ϭ�h��)���=l`K����;uK��]���>�~㶖�(���P�,��'T��q��^����T��ON=t���7z��9;�g��'�x�l��(�����j���ā��
��QS�y�P]��_�_���4#�a�٩��\��X �Q��" �j)�4��P²�ȇW�ν����'U]��� ��դ���B��,�����f�O6���p�W2�!��|^�¸��Dj�����*j7��#6|=��->ˋ� $-�\ Y���q,���P+PLW{�7ʄ��z��e�<]��b��	A���S6��eCAAy[R��M�`m>K��ז'�����E�(L]jf)�/�e�CS����>\��?L0������k�f6N\:�SE�3+H��2�k`�PG���0Eڥ��:�ԟzMm�۟�v3�����ﳲ��Wj����w�����=�E+�V&��֙1k�>V�!�O�)����Q��%K$��2�JB%}��+���,����[^�g̘,!��b�C��<�C�f�6��;̭i���~��k�ḙR��Y�Dm�;��B�/4y�Z��C89��w�H��i��L�D_��@u�&�*�O��f?��*��o"�|�7��S�x�� �	��=]Ni�등��uN4����͐.�[������3=x��PS#�?$����n-*kI_Q�>�0�k`�;��*0Ti��#��݀Л����qk�9��	!��%����z��3���/�n�^(Û�L��]���������r��-��j�q����a�!eɐx��X]Y)[�g�ou�h w�|�Do�G�\Åb��?ti����QpVf��p̱�/XM��<c\AN�@�`t�#5��Kpߪ����
_
%÷b�\��Rwx���k��ƺp�����P�yh�'���\��uT��^���UK��v�0Q��'��$�$�R�VTw�� Ë$�:�n�Ubɴޡ�u'¼] #�������#7�Q�@9��I�}PTV�+Q���1��MR�Z�Z���m��!*�!�	m���6i��Wx�2b��9O�J4-��Љgr?���%F��#|���Ĥ/S���n)��}�S�bie��5��-)�bSshf�,��������9���	LP��Z���
y.w�ӯP��i"T����2�e�P\���,h��;æҩ?^H�xmQ�hp���y�KQ�u�L�{8���r�G��E��s*�ŮL���\Q��Ѱ�̬N�B�SL�����\'G�G_y9��P n����i#���d��ʲ�#7��	�A+M)l�ل\��M�����~�������E84CS�|h4���&�.�A	sӋx��������Z;}�^���{;�'d��yl.Q�[˱M����4Z���Ȧ��~�ش���[���;��VJ��+�*�W�Or5���`U$��	�.���Nw�9����v���4��A���*>r�'u[�7�&�߃������VL�I�W��{�ˣ/o��L̆��3>"�D��W�b{s*�IΧ����P��8r0e�8��Y_(O0��)߸ �s�ى�O\��&�v&5^xYk��lr��  � �	�c,Hmms*.)��n�45D�d�^ʭ��v#�k��>�
Eɷ1ڕ��U����bN7T��w�%���д5�\���(����,Ć��Y�O���� �U2�c�S�?T�풹�S�cw�_[?1ߣ,�-j��:�/=.�R�����1ML��[�����0��*���PK��*�2ɥ�Ѻ�������	e�w�9���0�Jf��5�8�%{��u߀�PU=N���n��s���ڂ�DHJ���͌
�@�����6��L�@��S����)����_Y[��Km*[��Q� ���Mv��ϖ7�J��G��T��#��}9K�Ơ����~�믦��ʓ1T����T��c�B���Z�7*Y���1��0+�|U/� W�,p 8���w4F�M�cEF�^��HaH��:�3f�^E���q�����{�4����X���w��XF:�c�EC\a�i���AC���pJw��=(4i9��Zѣ���Bd �W=KȾ�r�ԢY��7�X�7���ė*�P%m'�#�0 b[h���1�a��e=7ZQZzZa�/œ�z��R=��Y���tgP՝�`�$��������}!]������6j����+��C[�}���r�jY�۶6�uTNN�{�� �����mM�*�G���ݶ�9G-
��x�0�ɤ�Ǻ;��S��5�]B���-((>��|A��7VȽ�z��&�%��;ۇ��撙_س����I�ꁛo�����d%�}/����k�K�M��S�`���그�A��t_m��Z�"S��x�/�� �����l9A�K]��s�Lzt��j�!���Ƅ)��<�W��5&�������'�2����v�ڽ��0���F��$���_�l��i������J;�J�J��a�3�j�1��Mg.�A��A�f&��d��ZT��J�F>`����e�0~�v����]����5��^������c���9�����"3ߧ ����{�C�ש������fM�D�Lg�{w�;���j��ې1�z"����?:Wt�����*)*7i23]�S�
#��U���T�"�[���[�r� C��!�0�x-�E'��X�v�&ff�h<"��1�ݻ��O�����L~{���\
j�w}���ƽ\�.�qsY�������p(��c*ll,�CS$(OR*��%��6����be�%˶����bI�.f�Qwz�}u[٢��As��N��j_.���g��#��Gä�@>����EEMH���?>^r5�
_g��<�=C<B�2��F��7�A��i�_]��E��e�<��Ϋ�1�3M+G����v֕h�����v���Kn�jA�؍\c���� �&􋃿�2$BC��pTQ���&[�i*����=��i_3�F8����b��TΈ����\�jI�ߘ�J\Xh)��_�ad-�iI.�~��Mͥ�2[��P�
4yPr,Ʌ�L�8=@a�#B]Î��*����������>�8�['��2����l���RЙ���ЕS�F�5��e󙂕Ŷ�A^�ˏ���+}Ӕ���/��:ԧ7)L�ɞǱ*�dn��}���Nഢ$���� ��K�7�Z@��)M�v�N1��_��W�D Ȑ ��!�;�_w�³�A��aZ���/I�j��R�Di�Ӡ���@����.�[)u��R��h��އ��Ak���V�V<���9��u["oX�D�P+}�P������b/����31�_�>bN��ZzRk7S��}�&w$�2�MpS�*ֹ�W��ʻ��"�AԶ�-D�MoR
���H��?�g.qܗ9~�-R�4S�����W�^�@�͹�2��1&�w�(ܑ���w�RYQ�����<2��A ��qu}]�4&��Mg�ە��2�n��-V�xy$�oR6x��v�gO1�RbE%�,R%I�j��e*�#�չ���4;͜�Z	�P5��/n�<=��.e�����Y�C�4'*O��c6ڒ�Z��]wN�5|Q���&�>�F��V	#����Y�E��_�:�V�w�8�Y�|#]�⺭Z�ũ�X{��.�ݟ����]�8v����4@�!˽��,�8lL�Kg� )r�c$j��+��[|o(AV-k��� wu"9�V�d�@�D���A]�&���LP�W�h�|s��f��]7/�xL�h��_�ՀR_��cA�©u�h�'�wc���X2��{���j���ܺLИO���^?��xwכ~j�`�%A���D�Ӕ��!۱o��F��D����)"�����?#!��
��]Gm�m� �ӰKݙKp �.�ݷ�v����ퟹ�w���U��H���q���fM3��G���J�]��?jJ�5of'���������>/5W��
�q�X��F������?؛���C�W/����&�ؘ�y�a�G�Zq5KH?�i:��Ɉ����(����8�g���������c.44�Й%�rʤmt�%4�ކ�C�^q'Z�D�[.�u�����"1�a�Yj`�湡2I ���;swD��M�2CtB�T}�c����\��c}fh�~��/�A٢�| !����a���1��}:���ҼV,�c�bm˗����;v5�?W^
~�=�-R���&�ljƆ2����n����V�Q1�}6�����N�GkA�P}{^u`��h(C^Un�N��Y}����1#�d}V,O2ԆK6=ℚ��*2��g��e�l��!"4�!���ev�-��ڕ�v�^֝��S�t)�����1���L��ǅ&&�p)޻��O��u����]�N�)�
g|g�Zvԗ��Q^Z��%�����\�/���y��&�;|jǹ�&��������`|�!Z�{6*Pޞo�6c��a�uyd/\,����R%4܇�/��&�5qז��Q4��3��j8%9�	�� �s�f���m�֜W��X��P����	���x������O���ea��t��r��q��HN8�z��Iy����QpܴiN���خaq��8�E����y����c�FI�E@�����l�q,��w'����O����y.�?��*���{|��wY������]�����`��\�Zy�0a�������	��@ �j�x������Ԋ��:�w��Q�p��g�mcGV�ۨq<��oܘ�e��p�����?�O�؉��~%�������M���j��,�� �ԛg!4ȱĐ�ˁZ�VؿU��Z��>�k}_�B�!��D�Kq� .������lP[o�H�3c���s4���Q�U�/��p ��/�z�-�շ�s«P�h%��CG�����步AF��䥻�&"��Q� �+���Yw�m�^Xſ-攢�Q螀��)��"��4�"�p|C��P��xz�7"��K+�j��ե�\���#)�3z~D�L����s�8��c�}L&��y��mю	(),+K�Z���X��m7�*�UaJ��#.���4�+Ov/�݊�Y�����m]�c@V����˛7E�fd�򓘻B����$g΀5����,n�����$8s�RކQ:Ek|�+s��+2f`�NGa�x����]�w~!Z0i��m<�VF~�$�-->V0�/t�������DD/l�w�b�o�Iv������nb\И��Q��(���T��;�gzA�s<�8�L�����h���»�>��0�zb�+�7��	�W1o[�_�c�j��ښ߾y����9E�QT�VG��yy���]dD���h����}������o-��G/e�ˀ)�% �L.�7��s��~ڲECv/�T�}Ց~�*%�BRr�?��{S!�2uDQ��N�H��LL&��ex'8��S�9�>(�2�װ�S�ù�-%w�M�����ԣ�AO�/�YT5�{�M���4m���߾p^^Rc��+���/M���+�'P�γ��-�r�+3�T?I_J��@]Ԕ�as����q���@h�4g�Q� L����{V�g�<�|q�>��l)�Y�e��ϋ�C��}����iA%x�k��Yk�l����b[D%(��!��5�$�F"�w��zW˶�{��JS˅lf"#��"�\P�<:�7��!pAߍ��t'�d�tg��G�d�W�(1'��I�H���Ԕ_r;��ăT���4�����u;N�r/-/q��wEL{`�(�p�X8�.<o���Q�+����Qv������!IJ���Fx-�b�:$)��(�t%и`��庹����<+M;�n�
�
�9��9��6� +(��Z����a��� G�xYx����|��r<�;��l��$��E�X�hy[$�\+Սl��� �j�N|_1��<Gq,2*-�0��1.+��5d�����Ӽz��C3e�]���▁��������|bs�����Q�0�M�|n���e�%t�,��-��R_'N�?���޾|S�=_S��t�B�������2ʊN�VS$����ʊo5�g'�}����vZU�L���P�����l(;> �Rs�{y'9�Z���&ץ�.��y�(�?4��)Q0�ْ�a��T� ��o�ı
�.�}�]�=�A�x�!�J�[��xyu��DK3q@ts������|3�щ���$��� γܰ�(55��G$�� O?�c��6��`�n�K�M���`�BxEֽ(k�)9=aW�K��J<��
]���� >=ByUEHM�XY(E�S����д�of��N_*�琲O�zѬ%(,q�3{y��&���D̽C��bk2�{�Yv͖�d�M������3��N�\ݭt��|�bHr�d���@�N��X[X=��YDG�<��$?�l>$M�?d�K� �`� U�e���]�0{Y�Ze�n����v<���@�2���,��&Gex?��[]�O�X6�S����{����ե'i�㌼���eܓ�(�:U��Wd�W  �!$+�T��t񙾇UTR����7Mc�ю��›cq7��3D�4�-?З��F��ELD��F��ذ�Yh")�c�o���Vi��� T��Cf�9>�8��0CW���7��9Z㥩j鋢���_]w����|�LN�O��v�ԝ�r�1*?Lo�?�Ր��ԓ�ƥn5b������*,Q��]qc+.�\N�V���Z6�I� �
���rROoJ]��g�g(��L�q2��s�9]���0шZ~6ܸz&XXI��/\h���.�]��xy�
��]�,��e�6�\�Eۯ���9{�R���x���t?���*{����>��W_/Z,�iZ2%����\�,��9�)o��ַb�@��,����$���"�����T�������y����mo�v�1Ϙ��5i��BYU];3��Ѡ\�~`rn��q\<컉���{q��-�����:j���C�+ �.Gʯ���<Og�	�r��j���9ݦE��g8�"�КIP���'�-!҇�FH���b��`�oe�U�x*I��A܎��I�����Ё�,��i�B�#Q�o|��-�4C~7�,R�A�]��e�?�U������)r�n�N��W���Uo�n>�� ���609��,�֫"ѝ�k�>��� �K炰R��>G ��B�u�>ubm��R��O��KѼ�<7d��ĵIu���n->�Z���o��jFe,9l�������G{�=��	^rr+|[��HL�u@!&�q�A�O}�:(^��`+J̓r��S�u#4�+�"�"�{��;��3�F�\&��Tn}�YV�ms	���:��À��m�J��NfpG�-���o-���E�M�QGp�B;zy�sJ�l�����fG����Az�!���K��8#F�^���
�>�����湜���nģ_�m�I4S�]E�R!j�qL3W��gߤ�}	�Z�[ny�*�1Kw�j�[48<��9�|�[r�Rj�y�H�4�q�~����^�i����C�XR),�����kC-��j�^�e����)�+t��:�wg�s~���ݳO	�L�0��
_}�~!\~!����M�l��9���-���ފ�e9��d�蟿���=�tj7ޮ(�Є,�%0!uO�£���j�X�\vu���%#��˼��	?M|�K��5��M��i����ul���>�7�6�҄
�$u�?Jv;�o����6G���5I
��}���l��3(��'� @�I �1kqhy���;$�R�]�tZ���R�{&���c��/�O�E�1/��� ��,�ͣk��Kk93!1����<Eiշ{�B�60?��*'�\PU�6��t6�<��vg��n�t����0Eȡ��2��I�|�c��h����@X�qP�-�rP�Ԥ�R/=������'�0�
l���VX��$��ƿуbg�r��9�36ȃy9qB�tR@r/�wmeǨ暖6ʧ3;�)�І�"�����'&�4���#K~K�2�#�������O�Z'e��0���}�I7��e������ȶP&_����՘�+��#��RFn�]��}�-c?�1��� wl�?����<n	|\Y���dtUpQ�k��5A��#.J�.��w�D
���E�{s+n9;N1$$x�qz0�,�Џ�8W�v\(�R�σN��p�Fd|QYk|���dN�U9�IYvi_E�0��F"h�ZEk���%���2=���g�Rv\��ғyw7� @�z��9��G��U�B:��eof���x��Q������إ?}�!e��oǰ7,c�������΂���i�}qrU�-����E�y����MoI�BZЩKg3���úF]�΢l����Eh<�t�-grU�A��У9n�\P��}M���2�!���6�XKCk���ah�����s�;�& �l�����<U�NӼpEڟ�l$"z��B��0�[5묇"������׏<Y������:T�4ao���<�+�a�Xۧ���V�B��w�%����%�4KsU��Q���\6?�r/ASJ��bxY��)Gۇvs!�@�虠�����瓈�%J��^})�L �C9�����|�CJ�"��L}BAk�ݻ��`�@�9��-ޝ&����`;Å�)�%[�>Ձұ$�~^E��1��Pת\~ ����zװ�hR8�����o2��j"�;�>��}�v���r3+���Vj ���[ʴ� m�\�1|'X�3�=�!fW�R�	��>��'��i)K��w��}钿+��;>���W\�r�,��k�.1uH�_m�Xc�@��B���'6�i\�9����7ѧ.�N�H֠�R:��Mq%��?��I��������'���;��lh�Ӹ����R ��������f��+@� ��nq[vN�g�����϶�����{Q��� �9Ic�i�*᱐����y�~�aU�S�:j�C��B���W�wk�n�V)0�m����G� ~��(E��W��O�)S��\�@��'}T1j�c�rS�4h���݈�_Ո�7�zyd+'?�A�GQ77���j��/�L�!MP<��ҏ�W����T=/GM(��Ǌ��:FO�bPk�ۉ~ɳ���{�9㗌c�L���2NG��ឯ��Š�r��l{��f{�R��62<��1S׿-�_��a������אm<T�ɸ�Nsoj��9�JÒ��OV��䤄�чRZ3#��˾{G9	���7m�T��"UU�u�|NoR+7�S��x��"�wn)
)�m���S���{{��H��J��Ic&�[l]ʇZ��}-�I��L<v��Ŕ�G	�������C���J58Gr"�Ӿ�KJ�GP(��Q�Xk����OEi]��ɏ�������?�Er��U��U���{Ʌ�D�'A�ffמ��4����õ�镛��S���*ؒB8i�]u��G/�hX��#vBJC�0�}\w��8Ƣ���?%v���/?u�q��ks����e�^\��S��Z��9��@(���	@�G�L�N\T�U����)Ngc����솳��i�}�����Q�����8	���"��<g�Pn�
�P�G�J��f����ȯ��0)��!&=νYИ����A�TDb'��JcŜѧ��MG7��a�N{U��I�W�ppp�/�5�W[�chm��u1�aHϥr���8�����a��'b��k�k������!C�I����[�\�k8q&�9�<N�G��z/ێ
����Ր���S�9ݞXJ[�)<|�F�g�?��炳�V�V'�օl��U����e	��,�t5��Y���Ծ���y���D���1���r�[�a7�v�â���>���&�?,�t>�i���q�7���j�8�n���W[��w8����*2�(	�=�������9yke��A=;G��$��3Ie�W��'8k<+�[�bF�TY��M���O��4�h���k
�n;%�G�㣆�|*ڌ؉f�}�YA�gf�X�N?�z��A����-�����s�c��Iҳ�l�$��{S�km�!!�n&>h��A�������Vtq����ǡ=%P3Zf���M���������S_�T!G7B��b��wEp���� z��#��7<��RD9-�e!��%�D�ۙ_c�r����K�߃��mF�a$rZ6�/K���0#�a��{� ��S����U:]�i�B�����6��� �]���f�Ȋ-��$~0#�l�\�|��n�Dx�bhC��d�)�aX��c�~��?���?=�q�6'����l�a����DJ�Nۆ�����b���;[�"-Pk��*`��A�TK_��y�A����::=�����)
�����o�W�/|S������?:;	t�"�D�]+%$�=����[�@�����~���dG[���dP�X��HT˛�u������GEb��:2;7�W@�a�|�!� �������i|V?��^�@�954����GS���
H{�l)�\�}T��wb���xYɡjU�l��N>��PA�i�C�u��>��ރ�%�r��kt�X+��%�uWz~/�6����-�����S��_²�u�D�y~D�= :Ǔ�*G��%� C��E��R�if��f��)�f`�� �Y��	��?<����
РS�6p'����:f	�x�pû�<D
.Y�?�-���t��h�{��c�����&�/)��Z�����ޒZ�> g��Q���*#uS��ӹ��Y��B��&�K�0$e+#j}<���"B/��	�Z?��p¤���ʐ�fF�!�*08ϏX?N_ү��1��G'�k�i
�䗴��Wt���EE�E;�&�E����Z�J�ZG���*R�7�7�O��[D��׋o�_��e"�]H�ݑ��X�n+�/l�ݺW��1�m�pa�m7�{L�mO��fԹc{?ڿ8��'��r�{�چF{�SCr9�V���`gѹ�7X!YIMUJ��Nc$,Z,Tz���EV;��DL��s�eV�(�1���եbHG̓�(��#X�����%��sk���q����""�!r�}���3d&�[��gwރ��{o�S���:���ɮ���M�h���+����Z����U`��`�hu,��� 'KI���R��P�`塭.������J��և��N�W �P2 ��d"Kz����nƲJ�Jf�����	���m�O��E���,c�,
�ÉY�VX�š�~[_T"�z���w���D��:	u<X4x�.M�����(SA9GJKN���5�b�ye#C����������߉��nRЖ9��-8L���S-��rE�K9	��Cr@� ᪔p�T��ǴöQѻ޻��=�u���:���\s}��%���h �y�TC)_KyE{\����Npm��LQM̰h�"�)�����d'/H�#�>.���oǧ���(�Iŷ�o���(*; QN=n�̱PI,��;���έ�R@]g���k�֠᭝������i�n���hj�h���(Ɇx��C��{jE,u�0�O�-K���W &��0fK���~����s�`0@�p�S�*>�Fv]�Q3��x�0t���R���
H�y{vV�Y�o���g�u����K�]H`{aX���.���ԯ�]_m��N*��*�ʋ	�9C2����a�N��iq2�rP��%��r�b�d�}Ŋ�û�|�?!��j�+y.��T�~�Ș/��&�����M�#P���=��-��P���<����z�$�Dꩲ�?��D^�kb밪��^D|@O�^S��,ʡ_��
P��`JU��!G�ra]��HFvGA�̝UWJ׭� ���h���;�ݝ�M������q�F�C�������mݔ�Z�5fU-���'7�Dl�� u�� 2A� ��Ň_�_A�]��cbG���(¯R��>���$9�� �70;�"+!B�f�ξ$��z�����|���#[�$�TC�X�H�TB���.Q_%����\��-�^��L����r���H�H��ĵ=#�������E�ؾ�~W����W��HJ[�"�P����7�c����X�K�կ�j�)��e�v�Ƅ���h<�mY�>��ֵf(��<B�b�pO��p�盔�J8\�|�����c��0�~��Qo�/H۟6�ZDs�u4�H�����9��L�Ff�T����TC'��$�x��> D��KAn	k̛��֗h�*W�yߢp'����<Iyj�l����Pc�i�w�픀3',-«�݄'��	:��b��?�Yp^d+�t�G��z�ȍ��^�[R�kq����`g��x�{Vv���e.P�_&g3b���i]'J� ��O�Y���	�����)�W��H�8���ɖk�ȾV�mL�x��=�|���b�E��}8���_���E'Ʌքt!Rs�D�B���<��-�?����=t�R�L���~H`m|��Y��IA��M˝>=!�(#ݣ�''�D�r��z廟��"a�-W��U�YS�vD��>	$+�֓� ��:�uz?���-{����M�#S�&^R��q�<��3�2���h={Qn`�Yd6� �|��m��ۣ���b��w �kǟ����:��s g硞����196���'��R���j�Q�X�h�[4!0�1.��2��������^^v�Tb��\�ׄ��U�Ebw�>tq�JeP���Ѷ����?U�ݽ=��w�KT����\�hV��fߟh�Z{)�J(���)��i��z�?�&ld����pJ��⩵�;����Ѓz��/B�x�����h~ًO�T6~/�����/R�uߪk���� ��ܞ�R������@�7�'��y�����a��Z'�0>�39&��?��2�|�O�ѡ3.#O����(Dh��o����r���{݆���7Y�ڪ2���&��9�rX�kYM^�C�:v����2��*}��ɪ.�|?���-N�Qe0kV)�*�{1��W�ᱺש���IwL=����5=��]�\Kq�c�U���ퟣ�g
.]�$�)���6M�'��	�
��2q�Pi���.��zԠ�`ƶ8���jl3��I\�c;mN��M��Iz�`���\�um�i���o8f)��X���L*����$wTaه$5�䛚���f�������@�B�Œ{���D�8�M�;@"c���߾���# 2|���8"�!���U6"d�m�[�͜�b�i)��pD�w�&��l�K1�6�;l�h&�#ک���7�J;���ie薛=l�#�kᢊ��|i�qkўP��y�?׍�zp����e00V����,J�l��U=���Ά�N�5{�$�e-u�-84�NTf�yэ7���?kL��tҧ~��X�����*��u��P����l=1�n�m�(X=hu�v{��s�I����?�3$;�JS��3Y�'*|����_n�B��8�L�^�u �j�����̸A9�>:�|Z;^=��q�z���qf�R��J�,@�\^f�}���~�ǲ��ٝ� |xIV#b�C�Pw*yu�}{���@�\f��2wQ�̸����������D�\���T}b'��}���X��x�ssα���e������[�5)��:������U:�����#8 �t��fPE��|�U�p�i>ǚ���������N�i6pS���>�q��O&����gðPqC���ii�3iw�Y?��}�l`���T�iT:��B����c";�L��N
6��2���<�5��k�ǒ���E���7
�_PM��I73G.�\ȧ�5%��������ᛕ��Y��e�oq��z˜\���ᷚ�a�f���[��胊Q������4��YR�����S0k�=vP���x���:�Z��I�¡��B4�I�I�qŶ8�皕#�!e�u�͊��Ph��(0󠳣EH�,�f������ڽ-���J����l�Eȹaaf������57�躣��+�)�,8��� �3ɪ���=���3u��i"�^�Y��ʻ1��O	���N����E�?�o�%B�*πQ+
Fj%d��T��N6fŃ*�z��i]Ő���n�Т�-�"���h[�(�w�c���-�=��=�*�sL��ed�����'͍׽�SC��u���Jý�{��S:J4�2����,��������!�`�暡Z��n�˞I"aT ��\�����ęvێ����f�Y���|1x0���V�"�?����;�&7-˒�]õ5@��ݾ��j����MSV֠IΚ-C�{di��١4�2�y�Ы$ރ6/Y/QP�7AM�vĝ�:�w�B�R�lkb1C�"��B8\�dG���E������+�w +W;�^EY�Ьt���/�cI�G�2[=�Gz:�� 2*��A�{�Cޤ� g��`���q�ՙ�d����s.J����!�$�e�S������d�W' ��kgy������v�:��Fi��ߏX���T�Ǒ�%cG�_j�\h�����(��1|k��1�`Ѳ����#���Ba�
}����ڟ��Uu�h&$8vy��x�Z��Ϥ�����2�S̈�������c^���r��w��	 �,h��5N+R1���>�X(;�]�g�ڞJ0����&���na���Q�m`U�nd���0���"�a7$g��c�8�M��D�ŅQ��&�v���6:�H/���3<�hq���~�N�k�Q�K��uVP�5�'^���M����9>f��a^�5��T���nF6NJ�ߺDs�Ȃd�$��O��}�� 7�{�Ie��.l�65Q�LٶU��(Q��_�F��I_'.o����JfG��r��``��nA���Eu��p����E�;���1�A��-��w;�n-=K�b�Ȳ������"�Y\��
�������n�V��:�b^3����<i��4@u?���JR��=^��m�=�,�h�L%�%ͷ7��T\kY �CN����\�
���4���jQ<ק�͈�|h�|�I.���p4%.�gC:lK�BJ��7V�5�o�,JӰ�3A 9�ʏ�X��~�cR�$a�Ԥ���T��?3��	�u@\�&�������U�p�t��J���5��f�P?�,�keb��=C����l0_7h��yG+�=z��9�>H�����ެ�������
^3~����lj���&H7¼��_|��vD�G���Ք��K��ad�B�)<���~����9ͅW���Y�b���_�Ou7�i��Gj�7p?�4��?�k��aZ�Hy����	��
�Y�i�um�;5)��WL�D�:'�s���=��o���U�����a�pf6NҾ��(_��[y<�0��`((�ء��\K�B��^F0����9��B�K�����VBf[���W�zyI�Rl���������m�T��w���S۳���FF��J�A�!�0b�y�?{⴩V��?5�1��6dh[Г������\AO#Y����U�;�-���q����CVX���S�Ī�C���g{ÍSŘ�`���ǃ�i'F$�L�΋>�$17�<(F`��:WU�ψ��ot��l����x�[H^_h�{ú.�H
�Q���(a[��6���Ӻ9kh.gh��ָʒּjdA��r\�(�Qʦ�6|d���^�m�Tl��1�(��`Z�p����6�zi��Zy<�F�>7h�Ȑ�(-�wlն؉��g�.���ǌ�� MQ'��)m��:�|��;@S��Q=�8���|Jf��s�A��;�߸��j9��y��#��6�jj������}��NL5�����C�"��]��7�j��E$u��$����;���')�Td3��^��R��xRm�V�����2�,�]^���ӈ�e�?��q�������0џo�y���zm��t�2���\Q�������\*���"��r	��W�ݕ̖���D�I��<�,����l��uR*�}F��7U��r�e��lM$�ic��t�Q/���&F�R����;j@�����t��I4�kx�q�0��q�|��NN�<%:}2��)e�����쮔!�S����K�����F�[�?F��q��}�	V%�y��d�%`3�Ŵ+;Om]ݥ?���Ë�����G&��c|+�sdt����M��f.iK��XU��uK�J��5з^3�s��]�{�E�/,�ɧIՖ�L~�J+`AG�<��r����(.�%�k�)�͌<�ͭ��ت�#e�Yoǣ$�7xer���7�'���*&틡~|�Ģ�i�K�l����nl�%�o]SD�&Γv�����a�uO�����S��d�%�1�Ű���5o�+���I�s��l�_G+�y5��Ø�/MiD�Ԉ�p�eN5*/�������b�6F4֮�,��[�e�4���|ӝk�)�a�IЍn{b{��4��ǿ*�O����05'�!\fET풣�u� �dlT�+�5&MF2���0YS�S�I�Q�s	�|4.21����p6�s���y���� �˗a8�y�e����2�`��-{:{��5}#��nf���Pe�s���YMai�=�	�U�rSHL��e���Zȟ��ɚG���K)��=��r��^����%��s�ўQH��:����`57nl<*eM����Z)i�y��G�g}j	2�H�l���Z�d[C]4bi;#-v��!*/�i���T���"��>g$�,#^z$����ŗx	b��9&��e�=Dȧ�����'���0��ݴ����^���P'jx��P���4bE`�����z[Zg��춬+�Ki��g�ԁ�@���xO����{��˯�V�uL24s���&,H�gtߠ��5�;|�����TѢp���Յ���Btr�p����е��w�>$����D����@��!�\�����w P��`Nw*W��)P�U� �&¦�6�8���_@��=�ղ1�&	+�ĹG����Ȗ7c�K�����|8�)�	����4�P��7x���-P������1�t�iwΊ�:�D�G�Ŗ��JH`�X%|�W�9V�w@���w?��w��'6Yqq�Ǫ���	wDJ,��zi̾��-ɹd��W-)%�M���X�
-����nA��g	�S���R���`�|�1���|��,�����w �A)�F�G��*�#?��מC��8e� <U�����PU�y�V��Sc?ʿ)���mp�٨C����[��l74���ۨu��U��T����r�H��.��_+�B5�b#r,刊|ށ��Rp�l֟�sE�|��"+(��x�,�W!�*q��L�"���6T�"����C\����_�qkY�]����^�۶��C��B�[�演�a]_⓾�,�JX�Ol�u�)RC�Hχu_�L�ZWB����'b�AG�����_�^OL��O�
��o¤Jͫ�kA�1�t�iS$@�E��s�5��__�G���!}�B�إץ��=mE�7h�g�(��ё�6�0��Y�%��u�ՄW�U�6�c�c뙏�	;�Ѿ�8Y�#M=Y��������i2��Vİ:LJ����/�F_Q��.�]�\��(��ϑK��VtM���a�}���Qҿ��r�SM��>�#l�3Oqkj�Z���vf&]��ŒF
� �2�u�(%E��5>C������D��n�;�����`�	F>�O�h����Q���X�(�>�j<[���h]���xX�c
�}��(��}�:��X���!��-�G��}���L%�"qw5��`���	R�ŵ�(�>5�s9���a�-\�?�f��;\)9���k��%�A�M)r�#�&����ܒť�<��56���:#��F��%��>�1Z
7S<<�F=�J�
*��.o���i��-�m�Y���� Ls�����qcä[��M��c8����V0��}�Q.H�%}��^v^�0�V!F˭ٚo8������7��+����s�_x>��I�j���y ���q��cJ{}�m4��lZW�l$U,��״���䡷�뷕�撫�Y��\*ش��k��@���F��e-6lJN,�m�WS�,�i��A�%�l�"�f����0����WN4�G�����1��٘��B܂G� ^��; $�%0��R����M�IU���IfD��13Q�� �2�ԎP.-���'�T��k ����^Eټ'x���{k��%�kT��`��,o��=�/��������J��A��+ة�W��	��LP��7�"�\�F�g�R%�������q+
	���ծ{�e�G*��W(8Ɗ!6Z�v��C�\c�TIBI� C�*�p8�����W�$?X���P�r*x �oH8�O�'S�&h�+	3\���>�㟺K������`�(�뾕�U]U۔�ь����g9D�@g��m�հ��������7	:I�M��v�%~�q(f�e#BĲ.�N���E�A�tz��Y59t�)Z�"vo�j�^�<������Т�'����t���ޒϮ�;�1 ��|>Xp|G��e���fɚ!	��4c*�<uľ �$�;�19Ow����d����r�^��:_���1�S�hD?�Y9e�N��.q!�h�N|�nd<��(�jѺW����^�,��A͗�^rp���M/>�A��%����'�8	�c5�{c��H�`9^�l�w@��-9�d�	HH ���ݬ����l~� [�
s|:/��#)�/<�q���[W~a�<b��cO�����4YcAe���<R.kC��	qLV����R���*;�;�6���i�;���y�	|0���$�c@�
b)��5�)}���p�=��rik�ꣿv�?�.�ۖK���ä�N�=�#�o��<�
d�쁾̊��FК����m+7V �/|��+�rt#w���oR�b�K��{s��p/�wj�%�b����ijC���
��r�QS��rj�f���H�Y��塨�W8MmOxR��y�/Զ i6�����>b��F<�O�vzd�%�а��LY<Μ���A�Y��|Ql�(���E*��,� >�ǒ(8�zx�l�=/�~E�c�ׁ�MS�!�*���<���p٠�6��{�t�O����R7�ث=�*�"g[A���׳zG�� �_<9�T{��)����fU-�t��NB��R�q_O�ի���JģnB^�*�������]�?cSʢ�'���X�Ü���c�5����߄����ď\���*F����=i��}M�����?8��uP0W4�F@�����{ÎBY��&�g��"�\^��`�_�.�=��B�N7d�<��?H�]�0�-��T��\Y��L���U��ւ�*�W
B�!7�MEk���s��Kc�e�B�9k��d�{��F��^G��h
 Jg�Ŝ�cE� ���Mc�w@Z��#�BW��/I����#�٢5������ߖ�s��_��esG�:r��p�	��R��z�u����̒�D/��^0���)�X�W�?��.�B�W7���@vK��V�Z_V-���z�rl���&"B�����v���.d���TL���7K�òI�B��* S8A�?�:==��)���Vɘ���mC[�q��1����FN�`��T�27y���o���Z�s�T&Ѩ�җ�)?f�}�~�>ql@4Q�.F�<~=�A.y���q�xZS���q����ׂ���[�ꥣ�u���JDIy�܇��9Y�D�-:�p�䕷������F.3$ܦ̺B"_,j��	��;�{��5`�g�s��pgD��E����K�e�%���xZˤg�Wuq���+�%o�}���1u
;Q��g���M[A�8��*ʄd�sZ�C��hfP����"�桲�t����3С꼻�z=U��x��9��u���R	_�!<T ����X��ixf��Q��w@������ F�)�gL-��!���<����)�n���1�C1�!�A����TPۙ�q�:�cx�~5,;�u�.:b�_�C�A���tZ��N6����>M^�
H;�;��|���� ��ʱkw��S�s�Zm�w��@tzl��4���]�sT���ɔ���K���7��>\���Xn��荜�rÃ�	��5c��Aoğ�=�:�Jl�[=ѵ<�T��ٹUנ���̤�=����BԱ����X'\P�XZ'$f^2 �B��ט���ț����٧�涎��g}ܖ�����e���6ʱ�݊���)��^Ww�w��j�����Z���M����bF�����
^��➵�%���+홄��g8��J�M�x�坞�]��\��p�-A2�Ř{���R(���_ q���-m�+��e� �������U~�g�'��Z�i2U1!��?n8��7����,	$���W?��!N�._��AՆw�%%���yő��(�%_��Ʌcp�i���v���fq�ެ��+@���s�θ[����؆:)��;uy�G��C`T̓�q�$�Z��S���U�f��[`�n�����~�B<k'U$�Ln��q4
u�K�Q��(w̽����L���N�-�dq��˧Qcwg��%{�XL7���cm���?��YO�5S��`�`�d����V�+l�����N�˽���BZBq��yD��m�@�dm�Rq���mD�_��W�_�u���9.����M�.�����$˷.�4���K]��_�| �S�9��*����ߑ��0����{rֻ'�f߲����d�����4S$VB8�c��y�o��.������l�<`���*���nkssds��Yi�R�|liI(o~l&��M��M �3Y���w`ɚXD+X�<�~ю35��0��f�(_=��p33%��5�-1�ӷ�~b	qր�Dl� F���/O���@�N�37IJC���VW�wVs���$Z4.d(�邊_�0��1�RWS�)�1y{�]i�sD���$���	v���H�<Q-��;����{�6wN��O�u_-���[�d�[��k�q	,,5^��ܪ#�a��W�6�S�DKI���7%�ƍ{^�Ⱦ���V�˘(��`c�A@A��6TC�+�!�hL���a�xɩ�[z��'���|g�펄i�=&���
��*��p�ه�YL���,��"��H9Y��oI����� �y��V��Ŭ�me�O��;��K�%t[���,�4h��l����c�Z_��]��4C��}��ss.F�	��"+x��Is��괣�o	ζS���	]:L����G�_Z�\e����b?�n�=I��Õ��n�"R�H��¾�n�84|=D_,D4L��z�~z}�lh��r)eQI��|z�
{�9,�|��I��m>V/�<5���
S����}�dM���N�`M��6��45U-Y�����+�!P4ZMbn�ˬ����w/���!�<�XL�6�ҧC�s	�~L�A�>�;�y�+�|�I�A�oS{6����1�Jl�t���<�3���� ��:y*mU�v�G�N�Q� A�����~q��=���߾��	��[l����u�2gV���O/���(��I��+�QP��xQ�v�~�V��݂������4Y�1�'_�/b��J���ʼ�N?ZI��2k�څ���xz�U��{�@ ���H�ni2p�,�y�<F&�/���6���LB�Mm�Џ���ܧLZ�����E�p��}�w���]���/��=�����Oj�e�����kS�����b�X�R��Q�q��J� .	�������65�6��(!�5���P8��*����_��X�߅E_��i���h���9f4w*������ҷ�� }8y�J�<#ɡ�ps�2�h[��idL��f<���ԑ�7�!�5v���=������ͯ�!"�ب��EoN�l�9����_��7󡫲B�\�ScX�>ԫ�#E�������x��껾��=��9���@����������5���#���ٰ)[�?�n���;�;�:[�Z�X�Ժ����U+힂[�����6T?��L�	}f�ԍ�D�x=�K����!*�oF�vv�W�Mt�$�q=a���agg=1�6�_\���>RE��\�Ȏ|~>�FLXa�����V��/P���BJ��v.�`T���.�J�W�S��d[�Ӊ�������I�?c ���(\~X�e���<�~tڧi��\�b̟���@���l�׍���Nqp?��Ɯb�L�M�$�Ee���YRHV;���K�j'~��-D?*'#� �f � � _*�N �*y�
o
1�"=ͬO�'w�7�sV�#�f�U���q}��>.6tU��n/�`�k��]���F�%mB���"('�<0�y'Oe�V�2JSEH���V��3����vup[� ��)7"�a���q%��w�'�U)�+�Q~��ِ�U����95X�.��XS&�n+��֌Ǘy�uր ��RE0��. ˬgx��x/>y��1�($1R��C>�4���IS^\a_�'�;e4���J\L8Ra�Վ�ck�9�pk7p���`�r��h+;s��܁��Z+����Rg)�(y�w'<LPa�ʭ$�<�c��uow7�?�<��;��h!���l��[�������90���Z�χ��f/˞w
.�/f?���b�Rp2��Ю,\3j�$3��l�ȹHץq�3���/U��~T����M	tR�f��9�u_�P��)u����
T������5����Wu�"h6]o������Z�wY�"�M)wq��j��SY��Ēa��&�%l%>,�<�4�q'<Y^X��%[z|$� ����'�UyN,�~Q�Z�6���ʬ�G׭�uK"�����@\��?��gS����zc�h�"��u�Z����|��2�i_�r@>�W�UQ�FR��\���y5F�:�������MU:�m9�>$B6����d�oޕ�?D��:Ԓ_�z�~��&��O�VI�ԑ�xbѳ��to��x��xU�Ի��y�L߸�֤�������W�V���{����Q/�r.�^������$��oi�J�L@��K���M��7��52)�����mq���;0�}"���N����f�-Ý~A�-+A[Õ(��֕i�~�wRa9�ȷ_5�ݎ/�ӭ?��{� p�ץ�]�_�_<ǉ9�(@������2�bw�bgG	��*���Qi�r�i(S55�S)�r�Ig����ƽV���t̽h�1�7��ϙ��mFl��Z��1H)���ȉǮ�  |�\P�§�OE����/���L#2���� E%W��w��ͱdq���H�8ҳ���������LaN8΢bᖜ4Z"5'B���zE��ē�Q��7_����K0j�sG�0G��}-g�ۥ�kk�M�M3�M��]�v�UO�����a�ؕG:x4��\e;��;�j�ge����x���f��$r:qzj�<&�?�|1��E�C|~��/:���p��.3d� T%̏�\��ބA��n�����AO���B�h�
����[���n!J[B�H�۳��M��o�1�դ`(�Xyh�0�.�E|7�������	��8�e�0՘k�/�_H9|��sKu�SE���E�I$t�yQQ`���g�ɷ	�K)�0�J�����\�,7���c��K�"�|����2��3pqnC|�?ΨQq/P�>Ww�*���[�y/�2V������vA�������_磡��;o�d09�:�O��&�Q�1s9��+����c���e#��gj��s����up� t����n�,��k�����̖����Y���5�**���5n�;���/se��x*Ӿ ���"�n�j����
�G�@VE;%��
���t
�����)x;Qx����W�O+���^��ħL֪�ѡ��?�_�!�'�y��?-d(����Y���#I��T߲"����02:����۾2�_��M��X-.h-�2p�I�������W�v���mYn~$f���zY�Qti�R�-H�/,Z�UZVc7��b���N#�!�O0f6k�-&[��g~�V���- �Zr�sv͈0(����B0a}�E��uK'����
<�6K�\H�U/��h��3����b�隻�I�NV�6�B1�����s�
3�2���n�M���n�}2w��t���~��g��_k&V�9<CЃ3Y)J!X�N��v���ɍb�|����S%��3��������o��3D�F����n�F���\�I��{0������F=�ĻeT�嶒�	C�~�~��Qk�;
�1�����K�=�E�U%�6�����[�U������W��+�8�j��'b���C�W�a��G����w��
�cv�!2�֦�%>�C�-�T�C�)ep�Qa���ƞ��i�Ӿ$@B�HPj��!�����h��#�
���j@�!�B�����h\��#f+o"òR�n���+�i��xYB��2ZNvI�ޣm3NDm8��[�B�ic-�M�v^ӯ&n�o%G��������0�t�&8�t��z&�����}wځ��+��,��w��%44b�	8�m_��.�Lg����ڵ�^�A���u`�
-h�s����F�n*?=?m���u5�
��B�.q\f2X��6KS�B2h�\�9b��Bqqo���f����?s!��h����1yd@��2��}�gj#�ߐG����h�������3(�Y)���5{���u2�5���'36�vV{,�ZM����)	\��1��4}}�TQ���]_G�����0(�����FE����u�W��\����[w��zZ[��`K��0U9?>{�jR�h92�n~X�D�!ho�����[b�)`�m֟|sk�\1`X|3���z+	��^�z��W��\�,��S���g0xj��=�S	�"@��g{_�d�4^�fuۇ�ɢ�?�>���g+�U,\�Z|���M�ETzW<�\��E�kL�?��@F�Gl5T�eC���t	ӷ"F�6��=�x�Uc���7�ӿsG� �ev@�
�L��1l�H�1'�4���KCџc���j����N��V��F��3��ߚe=G�e��	T�o�Z�����?����M����nn�ֳ��;8�ap0�Jc>��~Kn
�Qƪ�'�2�uq˛a���pF�� �ۄ�t�<�W���鏢���0���H��1{�� �x2�#��1�'T��Q�e�k�"HC��>���O�h���@P��!K�k��_P���Q�Xc���i� ������>.X�o{Fg�8�D(p�' L%IV.Ky4he�"��}4Hpo��%+Q�ջU��>���>l
Y�K��Q��-p�~����0�>�\Ų:+�}n��!����.G����|�
�:�7 ښ��:,%]��,�G+P���BQJ3מ�5����K��=�;�e�Y�:F�#��f���s�_���/��Pԡ�x�;�����n�(I�xK�N�	�k$�����#��\G4�~7�ɷkr?�����d�KM���Co�Y�;D-	����b����0�6�f'�J��RY�0j����348G-0D�{��vK~��i�-�PoE3&�uP���k�;	����TRSU̐� w͸��Wr��w@�; �R4����;-����r�������q�/�LC��6�����*�9KJ��z3(p��]�PN������]|6��s�f�)
9����?�[O�8�ޣ�r�Vz9UK�@�Z�>��B)� ���;�غD+�+���;?�w9 ��S��P������9RL���r�]�Ä����	��"N���_��3~�WR�_U�_}m�����}mmj=�nY�� %}���N���+�ޒ�C�%:�M���_�y�`K���l�Q�{���U�ޱ�鎗k.*��X��HŖj��V�g?��$Ӌ�x�q���0���T]�?��@t�pɷz`�:g���!k��"��1�*�(jK�o~�P��Fq�m����ӭ&~��˲�řT��E��й�9|~��q�����l����_\��������E��Q���w�\ϿR2�p|;�[+s�S�O����K1�`F��� �s̘�g��@i�;��5>�������47+�9�O�̜N
E��݆]�W)P�.�IK5�t���a{�v�,>nu�kP!H�
#4+>T�N?c �]K��Ur��}T�ב�έl���\��']u����Y��Sѯ�fy&�('�K!�bi�jZ=�B��.�G����	�;�`bx�:A���הM;�i="�]
ok�}����+%�O)�%"�qcߦ�4��8rr_I=^>�����/��әȗ���<�?�Lb��A�1����Q���3h �� �k�,�Yc��0TqH�r��������d����;Ċ����s���&}�bEn�*ʧ������^�m�賰��1|�������R��q׾17���%lf����T�/rp�ҹ������_Gr3��҉|̞��"�S�*X8��?�ݕ�a]M�q�F]��FI�;kv<T�*��/I��kO����i$Ѽ�<R.��Ų�d��E�jrs$}>xD�Sd�\�&��<o�����:}=O[�E2��Z�-+�����7�~hfJ(���-�\�k"�cɬ�˘|�|�P_�K�����$�s�A��?b��,�n#/t]�%��O\U�T��zWz���l�ǝ�瘻9��! ���e�P����OI���������WDE��@L� W�����Ef�-���3U!����M2�C� 8^�tqV�0��l>�ɬ.�^{��&����>�뵪��+�{�Q���D�=D���~hWQ�ZS�����s�0����z˖L�<�lzD��m�:��>��0��i�������;g��w�Ϧ������UU����2�ۙ�u���NH{������'�pjz����<�6<����M{��D�!e~F����z��I�A�+���a���aH��t��A^1��]Z�P94���ǯY���
�m�3t1R�}��8���͒��O�#ISըP��^���&N�d*k�I�
��	"�Dx�wRX�|��v <ޱ��R%������̭�y��P��E�Ѩ6����=}�����T�1?��_I���]���66t��oNl��pq���b��>���/���.=��-/��j��OY�:�5��!��Xdr\�1�l�)����ω��\!�T���|� ��х��{}�4*��?�T-萁�%�|~Թ�� �ا�ߗ������a�;20Ik�m�w�W���������@�D���몜�Z�-HgK�]w���@�Z��c��mY	1`V�4�ӓh�a�b70^DU��N�[;܇������������������τ��K)s��K�Cqբ;�#A���xF3ot��0��f��݇��j�y0C��$���� �� ����4ٽ��_qw���a˫;_O
��˅ǿ��K994�>�$Rm �yq\E%�h��Sd�; ��";�:m?a�f�$��le���$�ԇ'?���� �^�����S�V������E�uUnl���\f����my��v~z�����qҿ��k��D�"������x��v�a�\;�E%|��3T6k�iK�*	w������e�k�|�%[����b��g�%j��1����G9���y2�����3ƒ�ǫ��ݿ��H�U���������Z_�ORI����З38������*N8���v5bfp9�<^�����&�&�!*��Q9@���q���������fB4��=�0Bsz��qYnn-0�g|����Ϻ��fx��ݜilG�u��6��K��w��@Us���tZ����"��4�4�A����L�����ӓ��#�b��L��6;�x���ح�>��ϲ[��G��U�p�6?�R�mH_��[΁�L^���Hbg�7� C~�=�������Y�E�}xiEA��C�YB���f��\BB�S�v�����sI�^���y{Ǽ�c������5���Q��l*��3����b�O�G���V�n�詃�w��ZW:>���p[8��A����:��!Z�0��r;��aNO���89����A��=����w��u��t ��Dw}nź=�A�mn��M�����jUO���9�$�څ�&��2�f����ܿ���x��3��TE��n��х�ډ�3qw�iw�YA<��y^��q�WV�}A=^=ݯ;!ɫ�� �}���Tnt[�}~��n�L�5��>hDnz�ݒ�j9�'�������Sr�s�Xs/�.|�7�b��x�gb���B�m�k���)�3�����lz�c���8�?c�����/�F}�X(�²&1�jY�y�e�v�@�b��YefQ^�8��橝s�ԭ��!�VD����J�OB#G1	yq�ҙ����*s���.`F��-;e�;�JZ�JP� �D͆��$��X56���v��ί�$�����B�$��0���@��NN� ����.����<�ћ�Vґ�eb��'0{΀�9�F?�*�����I�S�򬏶���֛��+!�85w�dh8Ԯg2:�ܤ���~^��)9W�����t��?�f�] �o��RKL��c�~7�(�@a�9���X,�7�էv7jz�5AZ>�����S<���B���ݒ��it�(�c�R�Z[Ïc��?ϑ�i
�!s�m����.�N�\�������E�����t˂������b��?Y��ׯ}[�ϰ�0E~B5UAY=�|8��$�����3�'R�3ҽ�����>��c��L�siv"Rn�(�y(�E�!I��
 ����@N�'�CD�Κ�}
`(�EhgAu���U�R�C�|��Cy���lP���
ﯵ��6�<5xf�"6T�V" ��3��0�U�ou!��^9!Q�*L�ٛ�HC ���i�~3LYxu`s�#@R��W#��8��l�������8@���K�t"s��jX���J���
�C9��m��>���tgH����>3t��l]f�%���q⼷4ަ��w5^S.�zT�w�T-	��D�����y#a$]�l�@�N����q�f��g��h���٬�����_��%[��WW���+-���-6�:[��r��>�4�-_(e�"EgH1G�4,�W0%�|K���TC�8r/ 6��3vȠ���ȕ��uU4��;�.t�xԿ���v�֝Ņ�C�]������w�g�������,?bƁx�30+#�#^ ��Y��W�]
p��W��=�����d�\/LYw����eԴ���{~��ײ�C#�}]��8oF���~Q
�n�$;�R)�oA�<�8JI�,� >*V�J�!K	��v8$��~&ul}~��]�p�m~����Yv2�;����6vzr�z�,��3���+�GBY^I)ڕy<RW3^a6���h��p����S��b��˰�W.������l@���⌏�@�&�,��e�V��=����L�L�d��1���SߛJ��y��wZ�"��s�n33��?��C�U ���|�jm�^A&�|1�Eq��"��5uE�Ą�����:�3�*�)���\���P�,���6��w5�;&����E�k��B�O~d1!ݺpLR6YSE`Q����@�����O�����T%�/@��u�y�8�Qpus��"ʶQ�Է���+����Q�)T��K�|���Q��6����;8����5�E���}\
(����p�T��J0m�f�k c��; I&��&l�􏈟�k�C��w��Xj�(,������}*�n$	����=K-���+��{�!'ͧ�����я�;�94@��f����'�[�ŵ�Z�:������ɵ��B�s���T�Aw��S���<�A�5�>O��+n}�X8S33<\TY��m<��Fd7yM�����ܟ?}ǉ�$֡�����S	�~��6�?l�C���~�� �9㴘���ƀ��v�㧇}UT�/�f�sX�HX����F�)�?�x�N\_>�Xi'�SY���Ox��S�c~��*G���NJ�y�lb���T��@�㒢�ȱ�<�[���	�m�7�>X��j��ӗg���������s��	w΂Jȍ(�~��<��1�o��8]$���j$w�9���ET]`'��0�	\���QR�#�1�H �r5���Gf'�T�Kb�k��(r��ɍ���]�>z\Ss�Dx5�d���Sْ+^ub����㔤JҊC ��=]�|ZE,�/�:h W���F�ɤK��'~=?�A�52���G�XU70�,tm~�'����m�	��U�uX���M�_W�$,��)��f��vȌ(�Jo�����;�����_f
�I��E�~�MKs�`���:�`U��;�J"aB4JS����Q�(k��Lu�_CPz*���Vy�,u����d�Ah؉$�Ыt�,�kC����Z��(�O��'�<R��:i|�w��G����]|}A�!��$[��ċg��ű�c촇�#���	�/}z�?�B�k���[�o��ՙv��=,�����b(6�W�8���t�G���3Q�R{Cn<ޢ���s���*��g|����1>��^>	�GٻϬH�fT�~��/�@�\?�,�;b_���ap7b6C�!�Ŗá=e��F�!67F����Ai6?�3�S�_����C5xPS5�.{�ֈ3^Y[N(�5������࠹��uVC;�c�,m�'j,�o�X9�"�̮8n��;�`Az���j܅D����=�T�Y�06f8���'(ٰ�N~�V�4yT6j�U�:�.�J��
-;9�Z��c����6�����K���J&jS�.+NU���$>�.,Fvs>0u7j�%\��V6I�PTO��0X�Dr����=��0�?��|KW����!r�]��)�k�`m-7�,;IP�Vɲ8[��KYy����3�����t��5���>�=As<�<ox��d��2�	�	D,�l��=��N%�##����_�U�-�����>� ~��ޅ\�	%}��"1M�C�K��X�_)�˼�"���n~�̗s�ݫ@��:��Z;Z"��{a(��9M�$Y�g��U&Vcy�ʧ��fRM��LK�Aa�ߑ�E�|�����y�?aI��fS8�����D�w��<�M'�!��!u����=d���0���c��Ðwm���4
i>�7e�VY�����"z�ҥn��1���O���<b�К��d- ֛����?jy09�I�yYq-�ĉ²�<:�����W���%���a��e(�Ƥ��Ĳ?c�r�|m�>�cѢ#d���(䅼�ȉu�$`e�(v���Ր��P�z��qr@��]�����Y�#"���R4��������տ��M����q��[t���U���9�ׇ�=��/u�4�}vGE��'��mv����赜��ѻ��ܩ��O�c���5�M�!v"2��LJ^9��A��=gߕ@$�Ӳ&,sI1�z�b��	{�xR4�΍Y&��X=&N{��$�좂j:}��*Ŋ�D���T���dB�)-y�b�E����B*���I�4^v��x�8�[*������P�n��X}D X$#�����n�]�HQ���9�$��ˍA�NT�����U�� ��V��}vz`h04�����܌������p�@��E�A��D��t�|��/�w�S�s���O(-VE,���+�� �U�.Z��_�d),�W�<3
-�}ho}-�k���}�0{��q������"���P6ڕ*q�?If"�I�OLk�e�_V�w�B���CZ��6K���8]?#�^U�Mv-��moo��Ŏ�o�-�r)ё�C��|Mܬ�ӝ_#��Y����3I�b�R�*-�E�q}�Α����b�_9����
�@o���ʹ�VS�k��u��^����߸+h��c���t#Jv��d�W�q��9�ߕ�;��b0���3(on���{F�����3�ȡ�y����i���m�H3���k'�r��,z#t_B���AL�z�:.��߸	\t_Tp��>z��/-��M�Nt��+uC�J�v}�� �譠%O��i��bD�]MH�Xݵ����6R(��(��>f�P�&�2t�L�'�\��"V�!^7F���O��\�	>Ɲ�������c�n�ZTrfW�	(~��8��VoJk��E%� ʲ��Z�Y%�.&��z�bm��[�ܷʶleL�c!T����Z�����@�3!H�'�m���8�!��uǩ��9;��7�� ����-@��|���́Yy� >����Ν�0Ά��3O#/Ms��	QIFˏ�1d� ��6R�:&-�K��E�=�O����,����gF8��*�@��1r�>��3Q�Ў����u.��2�㹡�[��;���C�ɪQ�J�a"��n��PJ=s|����Ѓ�w� �1bwZ����"_藍�-E�!��C	��U�ɱ:��18&nD��� 9�'��X�#m�s�R1v{�]4đ���{B}�CYW+�X->C�[܏	
�;�J�����G��#�l�Pu��1C�͖5�87�;%�w�O�Ubjk�a��+��UE�W��W�ć�W���(��t�����J�,8�Л�����S�ȕ#��X�Z��T
�bˡt]*4a�X����Wߚv�:�BVqƞ���f7AC�ˑT�>��o�)�.���j=Nt2?v��������lu�.�7���G0�-И4���{3Ԫ���b��D�LCy�� �^`�C�<���&� +�?�8Y"�1,6�_�Ui���h��O8	�e�3�0A ��C'�fs?9�	��33�h=\h+��n9���u�՞�(���C!�^۱�j��6��=�)>EC�����$�U14��� ݀2{��G�6�[�{���0����j?Nd&��ɯ�2�jAb��p�DleL��po2v����۲��w٣S��S���l�g�� ��G�4�dAEkVƱ�CTp�~����ioJ��ɴa/��Z$)+�h�X:��^�>�cԷ�f�&��7pP����ב#D���������ˍ�F`����e-8����!��E�.�PW�|VX��h߅"ۂ_�Β�!��ϵ$/�<u��r�x>vco=�^��Q߾9$��]��T;���SN�$A��fu%�n����q`{���f�;�Bުpf=>��5W���݁��F��Ѭ�Nd_U��? 'aC���G�d|��e��	y5F�T�,��u�T�8Ƨ��B"y��r�wm̫άcX�K�m��o�nc���V�tWU
n�����]�/�L��>��QE�A5:^aCޚT�D
^6�S�bC�x���䷟/XBw��,��G�����c/�?���nLcz��"L���z���e�����T�ʊ��v�q��>���1�8OW��+�L�*)���/JY�9D^���m�%�x`��Ѹk�)���+b:����J���5��Be<�<�3#�HeFv8���>��j?���ǄA��c��{u3�'�]t2�_g���Q��wTI$=y��Fߌ�n���7a�QѦS�熳>a��3d��R�O��� �ӤңK���c��r-<�LF�R;m���SͲ����f�{_���bd$#	�r���f�J)\��t؆@�J�i����$H�zs�h�)U��;a7Y�����kW�"X�1|����t��P�`��=��w(�&)��6$��G���'�+��nu���~�t��v�8����E��Y^�A1G%���D{;��u�?�G�������p<t�ْn�/MB_�En�͔& �P,�����}��yR<>��B��$�4�t���� 瓧��s���ꂉ���rh�����	�����K'Ȃ=>Z��꫻Nɱ�=HݻU4]���hg
�����Q�;�J9pQU���ö��-���q�{��c��ٺ�z��|0CnK�ˆF��`���*��.+|���4Hw~��9n���޴�CY�ҍbcC�}�m�N4Jl�G��`������E��K�bf������7٦v������8�ڊ���H�4�-�^D�^�8S�+��?��7�F�u���/��*���������Bm�OJ\/�)��ԓ�]�͔�'�M�q֣bc+N���b3���:��xu������Z���ai���X�1�T����Fx��S�*Cݱ�q+�G��k
1��r���L*E��� GT�j4)�'�Z�4��*CU0=y�YWL�(�Ι�Ǿ�iv��WU�p���߼�lL��KUa)��MTdF6�S'kSYf�\�/�����R&�C�L�JqeË�p`6��/��t��_鮦,~��j 	5����v�.*+����Tg1��]��\
�dQ��է�2Pt���[��I��ϒ\}�����s������E1 ���?ϔ��MV��n<F��J�O�����O�n��+�zNDd�AI���(,_�w�)z�m^���*?`)�硣�u�v�#��g�j 6��_��ni����|t�J���� y'3���Z6G�&��kϭ�Sحj��b���}Qǁ|h]X���ͅ�3{8�o���W+�D��{N5R?��y�6�Ye����l�C��U��H��:�M��i]��O�X���&�W1�;;�}����b=S8�w���׏9�JO�t�Fӭ�����02����[V.�((���|�L�l����t���׭,B�9�͢��Լ���������W�	�.���y/꛽"|�@_RS�#�LK`���3�Ә�`�ճNx��
'���l�bpV۵	��jr��Ly�p�I��<f�P�������.�GM_K��f����u����in���ִ�n5��늏�-�׻
2RL�Hr���藶�߮���cN�1%�^bh�O+�.���^l�]!$��b �_�Z�o��(��Z��x��l��E��QD�����q��S$H���-h}p��d�������t<���9����5�X�{#��Y�=M����[FA�
��i���D߂���1h�o��Q�S���� q𮬖x��y{�,����*7�B�^�Bh<�6J�X���x�C,FȽ�$!Ž9��G��(ؚ}�j��gL�n��jS��MNխ��t=.�m툼o}�e��ie���}���r�x�Q��4؋�1N�9ʋ�X�MH.�ep\��n���K呥���@'dXv>��5���z3C��v H��s38�>�ʯ���������c��u�]����l��yұ�����r�q���Ĥ�M}�A!����5�r}�GL�@9,�T��g�\C ��>��Q��vo��FǖĉW�N�@ܜ*rQ�5�u^��^�[�� R�Mo�M\�O����{J�g,,S�6`�C�&+6Y����Qxb���ƺ	VS�(I������ U���`��	��h3\j
,��f�����0�*���Y�� ͞�Wt�$�k�?Z��"
�SS2B?���U�(1|-��F���o\f?�zr-xX<���*>�/�ŕg^Z�����	��'qy^���D��k3�9���z��mӉa˺�-?�=��2t`��D��T�6qj'��=��%i��$�|bD�Mz5`+=/��^�:QN�X�M�mڟ��kx�ޱ��d�6r�#m�cP~% �E�Kf2���*;>۽�Z������T��� �e_���z�� Ը@��K�61YV?M��ZJ� �KQ8����u:���ޔ(A�;ȷ���&E��+H�'#k��Zqb�z����m�]����{�G)채q5���,�(1�Wu�nίC$��U[���^��7(ɔ���OR�x����"�\���
��*��pxDs�Ĺ���Zb������ ���ٕ����V[.LWw��1��*��zK�yB��-Vl3���X�)�l�a;c;�'����bցK*��u�$��M��m'4��a��s?�㷬>^� 0aa��:%�;�_nu\�[/�|+��<�+�ƶϧ�f&b���n"^�����)q�^��a��e`)�C|q.KrR%��ښ��O���� 0�<�d����ҬLh���s�Ԉg��p}���r���m�vQ����|"kˎ���Ym�?e�x���Mқh���V����H%^>+��t,�o[[�yuC�	Ҍ�O�1��w�}$���/�7�i�ޭ�q1��4s~`��ΘrN�F�ez�\�TN�ȿ�M���_dv��#��7�xJ�xn������R�� f;����L�e������a�kDH�W� �z���'��޳�f���D���3>��jC�~��������Qa�����@9��L��N$ړ���pB���c���{���>�dh|��5_�77����$b�5�#�4n���m/���,>�I��1�c�uw�\ЎOW&z�xW$3�包�=��>���1l*Sߎ��A�yzÓ9,Q���͔�SHP���/:���ɳ��gM�>4 �צ?�o�*52���;��y{+xu^�:ځ�vVbA�~�p����xTw�i[If��E�%�ds��:�E y(�����@`ٓL1�#^}O����pH-�0*"��fY�5�+ 蠱j�5�;N�������6��(GH�x�o����2c�����,f�w�8�B�C�� ���jve�w�^� |nu�4z{T�UK���@�����c�-���.���}����/�R�w�x���,n_����L}�&M�5H��Gʦ��
 {y3	ꡕ�RJs�����a�����,B�n6V��p��Eh����B2���'V�lC��]�z�4�U5����+���M6�)��?�ψ#��E;s��i�j�Њ�nD���A�L`a�����#�3>ؤ�y>�˼��%�[��>��|_��'�,6?�CZ*Bu~L�?�`pl��/�������_(�@��⭪;;��)¢I�I�����c���f �6f�gm"5\�qyH@�Pʉ0��Y�(��ᔛ��st��y�~�v�2k��E�I�2�(I����ߙ�'���h�#]F���F5L����Y��6�BRߍz
+��)8�Jٰq8e_|o�Y'�m�[I�P�R�8��3K�����l�B`�}���IA@/��TU���E���{��Tq�I�ڏ��-�{��*/�܋���X��0`Q!�ayV�"K�μ<o�	D����&����]w.�����Ԯ�|-��E��١�n�=���K�ue�Ժ��xyȸ�|���Y�;V`1��z�?+����(@�����ϙ,�&���G�� .��6��<J/��jW*;`,��=�5�c���O�ߑ�kQ�շn��F;�$9�$ýr�sZo߂>L�vEl�)�!Ar�V)]�=�����`g�$�;�c!ߥlZ'G�I�|dH��/�\+�w�ֲ6G7I��H=׆m#��۳o�Roۡ�ZC���A�8݀���ڷ5���+:�zZ�_����XH���I�ϒ*��2�&
a��aa ����(��⫘��'{�>��!�E`�S������i8?�ã8�N"@S@���5����a6OKL@���[F��?��s��*�Ԉ� �@س��朄o�fNEDR��k���UK�-O��(��=�n��G��t\y�|�.~2JeZƍ3�������uG� _�#��t�#7��mz�O�/��y:�$��2Q�
��z�4$yb�}[X0�,��7eD���|��6\����[���R���
��$j}�wT��Z��{���kL��a��Q���ￅ��������o�){`���6=������VE�yV,�3q����IE��!����:���NM35��{l&��4CT.�%p� �Ԇ�����`I��H|�t���{L9eX�Y�8�����I���N��*U�x�V���.�egr)P����.���r��6���T�`�wJ�:,xY�}�3Vh���e��Z�E�q��`����w��I�O���=h[�l4�_ b?�jdpeW�/K�4%�}Y�SX�p�/��Z�l�3JV �8����Iu����G��Ƈǘ�/��,���2�,��j/� 3�"l�g,��c��L�W�_�R����D���>$x5}4Q�&4��m1�}F{�����`�47ILE���$=͉�)TĚ���M����?��f��Nv������^o���[��7}�[���yc�4���}wnz��-��M6���G���ϑeewOٙs�M j5�GB?�nAg�ボFI,\�"���"Y��� ��ge���$3�L�/"0cSx2dx ma��3��d��M������8E����?[�%�o��˃��,�#�s�� �վ���'��-��g��8~	���T
D��ƥ������:�Z��Z���>,�4��$To��w���ۨ6yA_ AO�'6��`{[�u��r�n��xK�p�0D��5F��>�oB�̩NKR�8�5����?Xj��E]���&*���Ǯ�D��ޱ������0�7��6F�,ô��,���z��g���µ�]oi]`������E��8s�A3y�����ٌ��]+\�������͎V�W�m���vB6y��{-��o��e�4����)�~�B攢�fW`̞���� �ܡ����X=�a���z��{��!���A��4��?[�jQN6�&�?B���Ԍ�����	1����	7�b{�˵& ���'���Ɗ�0-lv﯊{�'�e��=�&�Z(a�=Z�;ТE���S�sp�xNc�w�òU]B8�x��**���4iX�A�H����UK���C�lh{�d�jf%�
^�E�޷�I&T��]�k����)�?�۱4��hd�i��2L�^�"R�iiܾb}�y���ETG���it=�6A�@�JCF��X�a�����B3�Zl�k�)Z01.�U���M �H��M�ȶ� ���Ӫ�Ќv�_�5ܵ���6ӻ��a<3#�l��?�X��p+˱�,��kB�o��w�����q��9��]D��>�D9�f3A_{����Z��W"U4����-�7�,P�,�@q#%�?��YY�������'G�2��ax W�B!Bs�8�`�tg#%7�}���5W���8:
wk��Yy�2�&���B����d���I��~+W�aآV�&Z�K��9����Y�o�}�l�V~a�u�$����S���=3�0�H=��E�,l����k�-E�C-Q�rsz�r�&[�l�v���a��drΓI��Jh.�_��j�����OHH����y�L� �������}U,+�3��;�,F�P Ja|2��l1q��瘕tVw[��|��%*��T:·�H�Hm���*i����0G���q�Z�诃�� ��}�1U
9R
/�:��d.W�dn����q�[�r�B�F�o��*��!j�+�#�3ߥ��Y�߫�E~��l_ 
�\��=�s&l�S\6�|����b���U���ZZ���5\��I��.�6Fn���:']ܤ!�+��҃Yo��G�Sh�.Ʉ���	p�f�,N��m��ymi�?
>HJ���x�5v7+c1���tt������A;ЊX��d�������EP~hhDD������UBҨ�?�3ܵ�O�����"O9
���>nJ����wŨ�u^ۻ�i>�[q�U�U�VL�'(����L�����3ZjӴq�`�ɡu���z9g���!��f7�Y��ZÕ�a���Lĭ�nB	l������z�9C��'����NB�&zv�$�x��/��EXK�4�U�2
�d0�%7R{b���o�<�297�8˹�h��;S�kc��u��w/��[��V}c%�?�E�R������~�S*��ѧ��#�߃�t�Da�z.m�`}��u.��3����?�X-hȩm�-0��fxP��v��x��cU�}���T����d�v9VOWc���g�c(d��y �Ϝ~tc�ؠT�\�T�Ni����u|3�|��~g�,��E���;7�tR4,,	���m1��饜8��Y�d�SJr��5`��a����4��׾��R�}1�K��J�.�j?q��i�#{gd6��3٣1�f�>�=@'B��\3_�2��^�&��NZUoҐ�A�W���<Ws�&�Խ1�	x��d�ʒG�P�M���n:B@�rU2�-u����g���b$/ �S%;�L��m=�HHȦt��t�鐱�+9�"S��:�Z�ё�\�3�%�ǣ���d!���%�#V�8�'��G�W��\@	�J����ܷ�L�0�VV Bm۪CdP�9�١5ѐ%<����è	m;�9эe%d�r2���Kl�_bSl3���Xsq�;~�v�x�]����2l��=bX�0��Z��\��`��M�0��@�;��	���C��g "�Q��;CN����X���\x}�T��4m�e%��H�Pumc_����L�98�@k���}�VF���B���ї��@:��U��M������Q���4���ɻ�ӂ3y�`:hu�iYX��y/�.w�Lt�5��t��z���al�{	1+�{y���&�+*%2}�u˺�[q�"��#���S���"�f��a���Q��m�ϛfa+Q��'*�������ۅa-.X���C����z����%*�%!��m�x�����5DK�q���D����;�Q"��M��f����WQ�eju©|��o4�����	����/�����.<.�.Y�{t�ֹE_&w�ִ�D�Z��M�SsB�?UG�1s���$_���$����F���+@��Kt�wr����rEk��U��ΘN�	K��D����?7��d?䒤��M��+e_]����'���1{L���m�݅��\��XK�a�ԢUT�r�M�	�p��]��*���ܰ	y�B��!.��wY�����4ֺ��fH��(�ū�
�M��Ne��9 z�r���W���u�m�w��H*,�>{`��Uv��?��mv��ǳc}�B�It�	��z0�\F�S*b�i�g��L�.���
Nz/mx9�jka�P���j�hi#	Y�L[�+'�^��Õ�x���V�Y�B-!�A�������"յ� ��M
��h�e��$�����=�a����|ԅ��97�8 �5�� ��H_�O�c?_�s{-��tK�+��Ԟ>Je�%��H���љ�����Oj��'��;嘨h����-a���E�i����ۺ�@��4:�H��3�P�`��ZV:v㉱j���:����n`�����������)�����ZW�������7��ĤJI+}��ڜ�,l����r7�ˢ�.��
x�c7��]F��=9�\���|�1�����b&P/�%.����[Ṽ���U�r`�G�c4}#=$�8d����r!����sX���@����ׯ�m�님���ZM������v���4S�I<���V��m;w@��\8�+��β�{���Ja�k:,��%�hA�ۛh�!ن�/zo�x���G�c��2\ɹ�K>��5vL N��Ȣ����"� �_��#vb�ٗ��X�rh����#�
T�xݩ ��,���r�%�����ޖ�NFe��,W[�.�ܶ5Q�5��*w�2����M]Vү����"<Z�Z���O�1�̶�·Jo��P���D�&�5ޘ̜G�w��E�A"-n�,�P��9g��P$~ }|�٫yy�6���[�~8�!� E�>8�}���?�>���J�u	�5jx�'5�g�Wi�y?�>ץރ]��<�>&+~�d��y'�T+��M�*��>�핮c`h����{�vf'cR�e�I�� ���b��!����^����o%|�'����#�}��#)*I(�[^7>�NV?%mM�I��
EFi�.����/�23�C-bR�ր�����������s�<��R���Zj�cE��]�~�-�'�	s'uو� ����K/�<Q.��[+�E��%��'�p)���}�F�'�?-��ԭα�ED bkr3��%;/�q��S�³�/ CW��7�3):��ȶ��V:ݎD?H�E�F�|ݨ�]�x�B��3�B���wהnN'�+��p�Z70+���ķt?�(���D��lk��X{k�ӷ_覃�|������N&�
5��5t�*6���Z�L˷?��5��,���Ὗ(���O�0}{u�{uB'Rɮ%�Ivv]٭���N	 @���7�-�\����/G�C����FJ\�����^�{��{�Y�N+:����Mw���U���ƛ&�Z}����#�rp��!'�����,�PLW+w���X��E�%�l���?1�%��.+1H�.��c�L�OC�I|�O&�w�V��������}k�Ң��-59�=J�[�L���+Ol-5��@�=�A)+��`:!~�4Ŭ>�c�)��7JAӞ����V��=�5����m����p��2�xrw�o�`���~��V0"z���8hUyT7so�0o��fi�Y����'�Kl�f"t�]��fU�j�4 rQ)Ap1 t�nKy[>7\�������͋L�@s�	E�r�W�^�Bq���Nl�ꎍ��q�폡��c��6�9�ʂ�FJi���Bif�6�L6�P�]s7�(���C�5���%�T,����vэ.!���R�F9f���%n<<��5�>�2�ٟ�-F�Mgs��ޝ}1������~�oq�&�K&&!���-)��$�V$�[܈1�n]�L�~�a�4��P�E�f�r���j˷U���َ�a����Ei�Ѱ��?RP�3{t�_o���;�/�g$��Y���������Q��/>[�*W��g���W�B#y�mǧ��3T��,�ٲ�l~{�<�d�9U`c�7H@T�>w���7����v�ka�HQ���>�}x����"�}����̶;����W�V�U`FF���#�B��a-lݏ�u ]���.���4�v&�l��hV9�l�/�Փ3���y��ӡ,�������TC���?����f�t�|֘�=�
?����i�Dg<SwO����!��5�ɩu�����a���]� ;�O�P[o�����q�J�6�c�ՔS�����؅e��Ī����^�+2�
�P�g{]��.���2<1NnnT.;O��}h�����{N�Kj�J���{��+O���d�9��k�@r�PV*�=a�*�����zy��Yl��v��>������F�{��ށ������(�������wj/��(B=����O���ap���L���u���m�� U��-yU,e;�s�i�ڟ����e-��S����j����:]��Q{ѝ�D����M����03���H�a̾�z��H��QnL-w״Jt����Qw���Y��ٜ����Ņ���2��~�_J�=�戦?}��<��Q��i.�����1�H30��T_$� �m �D�@���?y��=��h8�4��kX��A�|=Q�;͊�_���x�}�Kg�+����9�5�ϲ��Ȑ8�௒��:�Ď2�� �B�GД��YBV�'�Ϊ�h�	��TZ��Og
�%���C	�Ff�{x�*W��%!��N%n+���d�5K� �m�_[G!��jJ���Wڦ��$��%)��_�X��g��x�PJ�j��X]㺗_ �^7��h� 8�c�&�??����J&!ވ�����hfԵ���] Y,a�7!fѰA�P��}ψ8^���W�����|�7|�%�j��$7?@���kC^i�m�$�\�rͽ�&�Į�\�_�C�~�v����#IpJږ�Y����+�s�:MDfo�s���L��dg��t,P�rsJW)M�Q(ε�'�\�g=��x���Qߛ�����+��[��h�"#�?y�v�a�F&����l�Do���-�����xW~��dcQ�O�jL��'�����d���@ġ�#���t��F���@��]:�����%��dF�(�*1����Ἇ��-ͬ%Jlq���F ������T|�5zy�.�!���^%�@�rN~$�s��c܍�YQ>䈃�Bl���F|I�@q�u9T�$?R���J$��n�b@��8yy$2�g,}u���oN�0��.ٿ<��M-I��N�Nm�IF���H\5֓��%���=��U�_=�O�^���=D�?澪)&�vp	���<�ww	.�]� �u� �����`����0��ު��y���{/�U�[��ҳ&���w�N<��^��`&��Ҡ��,�/��P�^�srK@�69M\���TŎ���-	��:���mb��h-���L�88bw���ǿs,���SZ�/>�U���b$軁��|�e"��l�����LM���p A��r�w&���Z���3����Ϫ�f0���c��9�V%�M�8���9��4¸*�Ì����,��4I�9���/���0<l��uW�7��%��˗������N����<eO3�=���y�7�������KҦ��J��r`�W�,��My2�_~jnK�QN�6���U����a>�SL=
�,o����`����G�H&}�k�7���#�����	ͱ3��q�e���&�͔�Om�?��4`ɡ����N��Q,r�މ=ڊ�HҔӈ3�J�>z�a���xYUE}Θ�X<h�{yD�R���.��/���������M;�!�:���e��������e�q,�/ļCj�M���х��MT�p몼`Ǌpm�[��<�ɺ�ָ`Y�MQ�a�V�h9��	�%E�����#7juyt� 򱴨�?y��_voj�Ŋ�<w�8��H��1�_�@_�����h��MKh�x��>���F'G��ǸB��)O�/H�,��Y�4�oe��Ƿ��UP�d`__��~��_~S)W����l���Pj�Zy	��Md�VH�� <�:���A��;��#���/�K?�{�2���v?��jK��]KK�'sy�OR�b�Y�O��Y���Vڝ3ZrY8���tF��9ςu�����^͜��K���^ݥG����D�Wd����vz:"wP&ft��Zws(����*���n����*J+\�נ
}d�9�zZ�m�8�,TR-CB͝r`o�9q��;M.W�����&��M8�UI0���x=���1��O���u�9�k�]���m��[�)����@�mk���ۺ���E�i�q^k�A	���Zt�B-��3<����Kߛ\�t;]�}��Aim���e�E�!�$_�������k~6��%��1�GQa9|f)�'�^DMn~�M?7��}h�~�.��4�|u�K�j$#M��ڕ�D��m����)�L�	�x��be�X^��Ꮁ��@	�7*� �8��_W���Em>��w\(����*{$b�m�W�,h����<��9��Ǟ���
�j~��^�Z���"B��W�^&�\ѡZ����k�&gB:A\h�</+�I�A~�(�I9j��X�*.��g�cG��-�X~�IO��j�s�طf[�c��2��H���Dn�����ĚKzY���nC��mi1�`��}�6�$Hq�&�.��F��|n�؇�WZ���>���H'�&���a���ƛ~-����.GN�}i�I�n�H'��KN��,s��)�-�8��fH���G��G���,��h�׬(����!��?������p���dc��<����{�Y��Ft&ֿM���0�#I�E×��k��������>. �M�Nn���w;���i}�i�ܯU*�	�ae^*K
��(9AN��g��r�4�]#Ԕ���FZߧ�r^�f�����y�����,J-�h3��H��Q�FZ�\�0��v��;}��־π��(_�u�'`s����ۚ�ᜃ�J{	bKW��+�Ng��i�^���Z�?�(j�h�hj
-�R�O$�[�]A����W�M螩-�~���匑D��5�^.\��^B8G(�ϣu>{���4D����,r}���!a�j�e��d����.�����2��K���X����SK���F�D�� ���$���S:sO��ʼX|�Y$`��������
AA��?��_��AN��j���K��sIy0�~��!j��o�#|�"x��B	�ퟤ���5�(�|�7��h�a��׾ր�HVR�8�j����.ބ@���:�@����/r�CD�#>{�P��{[{��ѧBN͑�Mg!�24j|���{�|��b�'��,6�ٚ,D=�����	���l����z��:����͎��K�BA|�AB.�;��RٲƵ�y�?Z�!�#��s `��)_�a���UeR����{��i2�-��.W><s�߭`�5l27�Q��v�ߤzR*���~�O�#������,�e]�;�Q�q>��Y�Yk	Y����!�����c5����OQ�'�`\��5G~��)�� ��>�n����H�0D�y��S�h ���Ǭ���'�`���Y���c6����Y%�������clv�%����<>&>�|�==tVH�l��zz�y���IuY�4���s���^ꬵw#Z��A��e�mï<˰�%�r1�XJ�.���hW|�e��,�YhZ5�.I���E�D���5#`���9N����!ϰ�z�ۊ{�ZH*>%���oo.����ռ����;ǿ��s��u���f�U�mם��Zg]�|�#�'��b�VM�� $�\��'�ޗN9y^�1�:=�:��3�@��1��ךM�ۗ���䩸�H�|��v�,�s�����ʟ�����/G��nz������E-�w_e��`�!FU���0˃k���dVI$$k��g��3�����6����t�*Lyde��MK&*w������9*�D���z�!9��#³� 	�~x�r�,g��<�����k e@ze���(��'�v�i����� xIk���O�9I�6�O:4ЀQ�Ϋg<MB\b$Ly���n�����	��G���_s��ž����J���	S̢�L[l`~yS���u�k�.���y�#��������}��ڍ3K��v
���<C�^CӲ�Z)����Iy�_�MАq�X��H���j�"�b3o~)�Ry��E`J�Ww����j�.��K���<��V</cC�\�-�׽NI/l�p�4�T��qWH7��i�dN���Z������Pf�I�	3�Ϊ�np4�]m_]$4�5��a����{�A-iO�;m/Q_�Q(Hg&R*G�Ct����D;�$|�"U�p��ۦ���ؼ��35(����̠r%����ΰi����O���h��t�~��}N%_n�����]8��AB��m�|������?A�)l� �����A��v�ku�e�AH�-�Q[ė*މ��9m>����$�Ttd2+U��X;D\x��Y��F~2k�����P�w�_{�h��:HVS�鋈��M ���q����O� 3r����{����:��p�#~T�{���rc�����H����W�z��'X-Ac�%�/ۚHM��ʿP}���Ez���\���'/V�Ɛ)k�C��uNT�}�z?��B\�ͽ],]��9+���Km^�٪���#�K����� ����ءcZ�\�c@����K����ο(��qܱ�v����ʭ��GI��7���l:�>�W44��/I.�Qٴ!糉�zfܚ������(Ɲ��^u�0��Z}�Дu?WIM����������hnTᓨ�� ��L�չb����m�VaV�K	3c�*�������`.� ����rˈ`�髂��@�z_�8���.�@�[���Ў{'�0'Y� �^e���/�oj��G��ޏ����4-�R|8VI�/�!w�P���n~Ûj�ȩ���6�D�_n�Mi��P�&���e�ˈf�i�k�#]�H�$������W#I�ӵ�B��h�Z������x^y8,k����8����N[\�9�V��wYwc:���2h�X?���D�{Ͷ��
��Om\��)42L&��_ua�F�&wL&B_j�-�����9*�����$D�ݠ;��g0}��nm�K��e�,�/g��� ��G�ű���Zͅ?lw����=���+���]�e���l�����I�m���!�8����풀��J���JC����X�'��'�D>c4`����.���*�I(� R�I��2�m��CL�� �ɯ��·����A*��I�L2���&�<�R(^�O���9�\�j�LD����k�V���[̖]mj@�DW��R�����&���x5��*h_�~��9��x3�|��&�s��b�˥�씢p4����t�\�$�!�N�O���b�$@�?'�x<�2����a�_h����){������B���_k�57ˈ~9�:�h��X̊�
�`+���1t����1q�=�I��^3��w�m�tՈ���pJ\�{f�����8��ϧ��k\fO�+ މ�����C�y�F�����K	B9���~�\��ÝDw���$�OV�p^�i�B���.ݷk9�+o���ȇVDzsrz=�Wic��Zyo�̯G/ڠ�4	�$Ɓ>6�v6�	&7=cN��IN�c�c��:C�2��,��?���D�{T:�
iC���HriG�BC:6>��|��јS��W��^u!@����	�d�̛n�ܾ�3N��y��d=��SAF�[yN���|6=��=��l»̀v�/�E�Sk�(�X�-��0�-�տ�/;=����-���!b���% ,�5&�6��#*�gu��fp�Y ����I���4��K#:I�p~�T`ǲ���;��2��G�SN"�p}���j=�ۯ��Ӯ�+Ƕ�G�.��e�B�J��Ҙ\Ø���_��H���?����ҏ� �עs$ɰ|9�v�Br�bz��3�,њ4FM��<'A7J�$�iX(���bND����р&ÌDg�!=��6�z�/�dbxDdA�y�t��pVo/��!���U�{E���Z��q��?2��[�$����e�������I�ё����\�	���_�w^-i�k_`j|�F��SD�������ho{[{v�=/�,
�1���͖��hoqK��d��FLU:~q������k��(e�5Xѡ��D<P��7��pq%WѺJR�*K8��N�e1�J��>�dV����
QM�H{{��ֱ^,�(���a���À�<dL�>9��VA����6����HG�Gk���:�O��J`�Du�� �-�S�:1��_9=��x����-t��ݑ����,?<��\3jH�kw�0M�B�j�`�3�H"?�9r�֮μao^ߗ.1���Ͼ/��h��J�v�u�)c폙м��N���T�^X^�Ʃ�m�>��#��$��{��#�u!-�-H��(�x%�7 wRy	���<��v�sp�Š�ǒj*r���x�p��nq(c��`�B�}���v���6O�ɮE��/����o���d�V4Jt��zN<\ˢ����]`�&���x��6,"���80&����Ah�4]�܁]�B"��H����o=�O�y��&!i��U5���W��B�U�X����f��G�VW^턦2�)V*󂠐gF��y�Q�.@L. ����	��v}m�'=�N�X���WĤ����Uq��#��;8�Xs���&�%��b7���s&j�D(�[ݮK�u�>�M
c�?aUQ���b�M۲N@c	,Ui&88�x��S����Fw4���,�?��^l/=��rtF6f��u�k��4��.�4�<GMz�|�o�1�ìbځ��z@���s�_wZ�h�hh�!E0Wڷ8.���(���(|(�8���_��{I&<[�,�Tx:�1�U��\&^���SB���n?�g>O��vܻ��v�}�-���ة��ϙ-�~5����{��8�vc���Ӊ�{����*Wva�N����ǥ���f��K	*%;u�������.��17��Y��,�G[a��E18�����!Qك�bt�o��S�Ӹ���!C,fW�o�W>��4u�?E���57,� ���l�o㹷�H@��$(ĕ"��V���d+�7߻F����<]���g��w@�|�é��7j{�/������]�i�.AޘV��GJ�9ۊV���?���2H�cBc���7>٠�,�|;Z�e�o]Քӧ�Ȇ[����Z?D��|���Z�3�t��B$��kq�n$�gU�-�������_�)?�?�����>4�zT�8S<7]�p�Y��_�i?iI_�	��ܳ��x��i���4
��v�y�*�!&��ðG��	|�lBN#S�OzNYǬL���p�iў̛XC�����j,��cf���r�E��o�	�?�9�z�y�;���;�ܦ�y<g�7U���ȝ�/|2���8��!xũ���TJ�+��l�2�_��b�5�ع� �>0��%�q$�Yڽ}�F��D��OOZ���ݿ�!n<����*���I���8��D��5���D<{�k9��݆��K��I�JW�;�q�����cO�5i����c�� 1��^b�E���]m:���@M`���׍ְy�'m��3��I�Ry�Z�|�T�������/�>�	���jhY=�b��Z�F�>�ϫ����@	��ӴI��b�X"�Fڅ�o�F���ˑ��)v˪�|��0r�mW�&2Ξ$�c0���3UIF"��in�"��~sڼ*c�^���a;�8�!3'�fK������Z~%A���`�MCÀ������+�3�91�*�?��S���A��Z��^�k��Zr¦�� \�>�9��F�	el�`��@]�7b�܌��[p�M�yݸxF(��#܏%�`v���R�Y��-�q�����\�s��ma�5�Ħ����b��|h��	nLEQ�$�ş�B0�8����!��7�������X!-P�ΏX�vuϯ�V�`e���f�!�*��H<���~۞H�?��V8��������̠y♴���z_�? ��#��*ˢF��*�����+�zZ�-�C�s2A1���j����ȑX�C�֬���hO��w^�.���=(��PⓎ���zJ|ٛb�}��r+b[��PՅ���l-v�A�\�GJ��C[]�(�������_
�a��o1wk��e���Nv�r4G�W$0�m���P�a���i��X��z�*<��{��M�rI���E:Á��co����}�,vjxs˫�t!�җ^��I�����s��
Dl��*�� �JY�2_��'�����쭗��n�D(���X,�W�Pg9��`x�h���~�8���#�%g#Զ�4}����IV�h���yKZ��׾��@�����R�f��yX�{	�bk]��^{�t!���u��D�kf��D�G
W��aT���#�G��yE�<$�b����{��͡����݃6���d��jOރ��h�>�̰��ÙG5�d'��2��B��Y"1�$u��x�ԗ�A���j���Y�<d1Ab���w��	S.��c GoYg|��r"ؙ�<9�R5	ro3�Y3�|}�0�z�QCR�l�stZlI:s����I�J��O�3R
o�P�&O�}��`�}�B�u�p�,�_�;�e��Z_T[!���#&i@z�q�"b�\��� ��p5X����ӡ����\+k�E�챉j�@�"�j��qsw��S�����G�jgz��'K�����1i���@�ْ��1����;�������(�|'�}�o!nmF�J)ޏ�Yͼ;/*��]Ҋz�?�W��i߰*<sX��p^(DA7b�MM	�=!!vbӐ��u�w@r�����Hyi4���{1� �#���nk�r�=3�,+Ч0L�*�Ə/�*Ͻ�A!Y��3(��&�*]�Ǥ&�Y���2(9B(��?w.�
В��EF������ҥ����
̹�?���ʄy�*>��kć���=�Sn7��Hg3����Nc��&ʊ���Ԏd�hS�u�~�ɲe����F��i�=��,���t�d��me��;�Q��DT G��4�5��|�N>�Mo��}�J?2!b����G��P���.3#��%�5��֢3F���	��v��~ �(������ c�:L�0S�3�>��9��o+�D;��I�c5��d�?<�5�5Gv���8{]�y���N��[�F %����s�v�������}�E�*�9����������L��3��t���B���E�/�%�T㶜P�ߣ���+�i�`|�Q�cJ���{���N��J�oUER�#�򛟟�&q������a�<n�����
���sj;�]�dK泶��(�h��wv�6H�-�H�L�zV&7nҾX�Eh���_!Hn��T4���8�G��[F��V�4�ٮ����Ir���k7���-�0Q1a�03��T��3�="8G�~y2���3�3EN�S��	"�Σ�~��<�S9e���*��!k٪=D=R��1���an���JL�O]Ĳ�sHW�����m�/�� 
�gzɪ�B�=�s?��o��%�l�:ݍ-�3I���]JK������j�$to�)~ld��y��6I�Gw;�"�U�7$zmӀ�J��i��N��M'4B����Auϐ�<v>��BS,��0�zC��Y�x�������r�@����������8�XK.3��;[K��_����/���#q�ۅ\ػ���$�?�XZ�i�#�J�ӫbe4\���\��+��~+
��%	H�3a�%�MT�o�k����1ெ�/���	�i�"������{�-�t����{k��f�"	��Q_����r2�>�0�-����������_��8�,�>c��� �1WU_�[Z�����V�$UQ��j�E	��'�?���Ɂ�(Ǜ14�r�b�9"�q �����gGM���v ���i)B{n���љ����E��؁W� ȯ�}������g;��Z)93��h��\Ѿ�� �bޓ��C�;�����z����&��(��d�З}4?���{�Fzp!ut)#�.ߧ\vM��k�+���+k�3�ge-�da?u��fsW~��D��w�,Z۪-�'ty�W����Q�6�J;��:E�!�7,O����mP\
n&֫fs��+i�v4վ�h�N�݈�A;p��OX��|x���*nj�Si�S����@���l�����+h�	�?`ӭ��������G%��(�RF�}H�
e�$/���]���Q�B1���tCԮM�M��LOю�O�x^z`׋[9:�s�JM�/��6�㝥-`d#��vG#2�m�I������>�(
�XZ�o�}����Զ�PwO^�\����q�B��~'��)�MO@i�jx$���I;���?,7n��Q�׾<<vvzQ1�q>5i���珬<c�g#	�Y�Kè^��N�RI�)'m[a�q�qGFP��w@�\@�PCDHb�1��Y2���Tt%q?q���`˭'���[�JjȇRJ�T�X����>H߮��#�?T#����8�U��IGQ���=��I�H�9v:g[d�\�u���)�>Af&&40̛���&�\�~����szV�1
d ��^�@[�6eB�`'f���S��G�!����v�|ud� ��lA�w�%bl��2�z%%\/Y�#��e�w��j��Ӂ�/E.S�V�#�DP�!{��2f��x�h��͇��$��6��#�����Z��:5�4�t��f�*G	��t�f8���R����=@N��/�iݻ�������D��:9��:��s*U~B^!Oa%��K��,p��	@�A^�Nj��5洇�������;۬[ń=t�%��"6D�h��ے��U�)����z'4��wX�@�ؔ�����X��F<�rD�8�F�����l��<:h���"_�a�T􁿭����C?`���ѻ�u̬dyedOn��=; j��]�;�����Fc����	C��C�A<aE�&�i���z�R��uƜ��O�3#�qڄ)m��Ұ�&s9�3�{#:�n?j#��=�0W��W�8<���*0��p����K�����qq��>��*�z�>T�����H����A��˃�7\�������c��]��%f���sGI#A}\�������u�ܚ�1�Ƣ�H���I��#�o����Ǉ�_-ݠ�sN�Ԍ�b��ڡ��%�_���~}�H����?kF�ij}P�iHʯ�+�C5'�%Iμ�>F�]eq���!4�X�_�pd%sk��~�p��cu�+���������\ǅ	�K��"M��>$XS���Gn�%�Nԩ]1�V�4t�Lw�6 V/�d��������#�ʡ:FL^�i�2N�Z��V�����a5v00���]�E��k�P�6�q��3wu.���d�(����Nc��&�ڃ�Y�����_�'����P�w�(T��9L\6�c����Ӷ��@�HL@ �4�9zL�L(���5�P��0#$�渞:�Nڕ��è���i�>���(�[��}�6�q�7��ZF��A"�j���Gw	�J\Bįr��.�s����E����|���םڼ�և�<����:�y���g!�,����U�4قw �k�P{&A��:��(�BP)�� "�G�Bޱ! �QX�k�R%�D�Q/����<�V�~�$dm�==��V
��/wFZ_�dC�7�w"��3���
����q�犨 �ʭ�2���C��Va��45�f��j3Q�J�=��_���+�k��@?��%�G��u6��~% <�9뀿	�+7�=��K�3�⫀m���^��˃k������+����U;�i+#��딊��W,BV��w�$���� (��9!{���)�jVY��=�i��K)3O�z����K���s�T)@��6����j�)�?�l��O%�To���!��X���0 Ƣm�MТ?3O��M�/(��Zg��h-�	_"4y��&øI�T�c3��h�&EU�{=��%}8�n�ǩ��΅�������.���̀�[���*�۱���R$^�TE �<�B�bY����gY�^��3w�[� v���4�Z���ԤG��t�zU1�� ���1S�Vm^���t\�3ƽ�3��]���5�C3�Ql�� ����; "��*�?W����Yxn��0��9��V?���l>�����Զ��}k,@uє����2��|u|̳����o���/R��U��B��?+A�o-�l����wc	3ϣc���:ڞՔ��y���i9y�{�@L�WH�>���.ںf[�CR���`��v��~L1�S4����<���A�TW���$����d�Ap%r�,<����\�p{����e�&g��: ���/1R��DϽ` 'V�E|�|gX;��; ��'}�p ��mӋIi�����%M��k�&^��
+�|*o�ŧ�������a���Xh�k��)��|׀Z�K|e<M�>���;�w ��oO��e�+�`��EB٩�G&G��y���4�y�H����T�ǥ �X���!�Ԥ>:�����(}�s�w��y�G}B�����+|߼j�<rW�
ĭw�;I4�
\>&�q<�0K0�Qc3� �g�D-�����2כc�5�=��h��[�tM��3kL���8��6=z6�?T� ��h����TT���W��ȴ�%�ѥ �K�'���$��t"�R�U�0xL͂��n��}�-����0������19�O�+A��8�֛!�x�QR��Έ!N��W��di��E���Z\��æ9N!�+�"�1EYZ�hP`d�l3\ [̍Q��+�;1x��T�k����^Q#�,q]���S���@�}�����t��q|~���&�ZY,�Y�����։���״uvq��R�>&V}�F҇H��h	�-5��Z#ǇJ�Hq�cl�
�O��7��G��[��9z+I��*��q�qB���T�"ʑӨD㡱bfw����6����Z�Oz*�Ύ:��XΧRӅJ�R]���,?g����ab���D����,�y��
|i9�A����Жi��e�)�i��m��G�;���٘[�O��/�ɧ'����v`e-UG��z>�B3�P���g�~��ΗB����$HL�H��Z��R\�����Z�,BàziШ�t�_�T��4LZ�:�m�3�=�}�G��ZgKXi������މ���f�jf�E�j��S�z�g;>3����~�U	��Zh�k�s�����%�����0PM�QnLz@��yJ�0!����+��l��Lz$&�0�j#m�a�ĺ5�`w�M]���%O1� *����{�4��1�e��.��F:�qG>���<K㭘WN�7nӯ��O�n��v*�ϴ'�� J����"����2��&�<�W�{m�6�N��jm
�>N��^Z���������&\(,������~;�,��<�PTc�Hݍ)No���m��xdc{ʍ�}l�7���y���R<
ڍcUQY>��Ȑ	Z��z�����"�������ü{'b-�\&��׻�>����3��^}a���/A�������?�8
����TFˬIϕN�ޅ�C��D
�]h�|7��[n3�k0���D�f���MY�NTԋ|�l��5���#�c��nh�{c6������]To��Tΰ�cD�h�*��x���-E��̦VO;�-.L�2�s �.
)���n������(���}TA����Q�C��`^W�v	ʁ�$,y�x�bPxX5V��[y鯍P�ڵ1_�������;����1�����x��t������dɰìn:1W���ۉO�F
�����Qn��>���t����	ۖ��,�2�k���Iu��ی���g�u���ݬY|�) >�&�B�Yc�W�|b]���9��q�ެ�2���?�-�m��Bȁ2R�nj=��YmW)�dx�W]7
B]�|}�k�G�2-�g3��fZf��A�gό����^�����n$8^A�Q�[�ᥡ�I���;U#���Mm���rZq��]o����|�k3�s��)x����V�v-����#��syn�O��ҙ������?�� �J�O�b�QY��f���W�8���?2�1��3���������I��6�V]�_�=V[�[Cc���0��y	L4�~�Uc1y�\@,(���bg}�J���yLq~{�|��vA�(�Ͽ�\����}+{��5[%�^�!����u �@�� U8J�K���S3(��{��{�4��pN�@�S˗Ӂ$�ӗ�#� ����W����~��lz��3�'�bd��TT��މ���~���G�q��ӄ�e�[�l�����v7�^�f���b���M�׉l�c����ɴ�ʖ����.��NJ#r�E�xsݟ2h:��]# I����G#rpĎ��1�W�h+^+�q��Qp(��s�B�_�_{"3�Nf��`TOr5J
��7�ҒNd�+�81��n�.Y�"���^�Co��~��ʺ
�H����V%�J�ek뼃�i�ݙ�ɊD��d���O�-W�CQ�K����4�ܒ����31���~⭍��]ֶ����4M���s,��s�N���S��;7�∃�x���V	�*� ��z�c���\��Ǔ5'�]�@�1�g� j��"�~��)]��r�j2���)2n.u��6K��U��V�6 3H�(��?��Ͷq�n�C��m���]C��fI�/54�"�`.�$i��d��g��N�τ¨+�
#'�P�Ҟ�o�on��5Z~n&��"�����^���陸�ٓ��)�y��\�4��kI��ď7�]�W�V�o��'*.�~qBs��*���A}�'��E�s�׋�]Ӥ�RJ�m�l��^�����
��HP������ʌ�a�o������*��{����HM��w@��[B�?u���<��C�!X�D�;`��L�ON=���(c��)��%�JR��� :B�&gy��X�Uq,Cm�e�'�ƤALO�}�ے��j8K*g�+��Οm�����W�Ļ秳x�?�_Ō��Rp�}�BO�b2���lL~�,TIC�=�d�:�}��j��W�	U�,֡����5�0~�3�*}i4���3��P_���wv�>&}t�;����ڐ-��}�m�JLs����i�����s��7�Ut�-F\o}
�ps-/��/�GA���L~HDo�f���e1�����،Q�َq�����b!�(�.U�,v�S�*�I���;���ڗ�y�C:�:瓁�y�#�zh���x�<_�V��sC\�;��]/\擯�oU/����?,_T�7k���+�=)�(!3��JpI�hW�; [��b$�+_(I1�:�f���glh�`�ؖ��{9\Kl�v$�<e6�H�Ky�|O`���}y3d��d�X�������L�*�*`V�"��"@D��b��|����
#�K���t{�\M�]o��Z>�Q���@�'Y����'���	�K�������9|����U��ú����2z��rDӁ�v~�n	1� q���;���HA��"�d�ǹ����=�룯�f��컖��5��|#l�"�!�Z� ��w�1�zVzF�n�Υ�6D-O�(e�����J)~�!wVvDsd���[/��s����12���#o��7#َ��� 3:I�%��	��X���MϘ�HD$ڄ���x����E��!���I�ʬ�I�X��@�C"�߂��͡D�
,����A*��z���T���/V<H+#��t�����A�r�<��R9I�e��u*�Y �S+		_���Ƹ�t_��늣���*E���H����"��*j���&��V�m4M&�>'�:v���*�R~�����%�Q:�Z��X�h�қ���b�T ���������+|��3�ʪ&���UBI���.WGLȵ��AU{3�Vpǖ4$��@���\�� T���8G�s���Fx(� \ş�/4��AB=H�uw�c!��ҋ�L5�m�^� V%�[�RO����,���!yдG2�sE��������z��� J;=]�}�('�?�6���H�ͦ:}$�Ȃ�/Y��-!�״���!�e&c9�N+s�v���O�M��v1FG%ƽN�ӟϓ��Z�J)]^%9���3RiPI�Jq�)�m����ß^c�lS>�A�B�~�%��+��� |�J��	�����r����Ed�]<�O
Q��n$��9A��З}N�I΃���@�6>!T���H�!!���J��~$[��Q)�$��T�%����7Z� }��-�`�»P`��K*�/zN�ť�=h��R��H�#����V�Eg��H79Bi���j�
��\	�1���M���nm*��e��P��tLq�W�ߢ��u��?%y� ��Ւ�p�3ШR�U�r��B��7v�d]�kP�$y 6�݄H�ޛ;��M�Ś#�6Jf�7�c�Pl�sNqo�5��)�*-h#h ��L��I	M�J:�{�Q�u������?��y����l?6XH���	�7YU�~���}��̤�ur�IB:ڽ���@����F;�~�^P��C;��?����^6��gf�pn��ѕc�J),ރ�B�y�*${ź���?�����Av,_�)OF��sQEs��΋�Th۸r�܎|���n�t���T���9�6G�Q���w�+r���c��k��.�TU����˂����=�H�V����N���(cG�~�k��9�u|�V� Rv��?����4WT6\��s��&��<s ��ѱ��%_W�4����*��zj�ܼ`�Df.�}���"��߷십$$I�����r�8w��
����xjg�V0{��;��c�0�$��V��5kPtQ�����x�|���U'��m}�X02�K�̻�$�1	�G�J���V��]G������&��T�"DWjs���3�f�������tr����+Է��PJ�l�=l,Ȟ�ě���%f�����{�=��q��WV�E�ڠ;�{�[���Z��2�[?�w�*T��s۞����}��)O�-z����1����g���G���2O|T�j~�Gu�V���u����9�1�h���d��>�W
���`@*��H&��m�	{��m�%Q��$�WKDv2�����t+}Dr�.�$�F���
.�\���>ފ`gb㜘*"7\����|ju01��	�W-�0��80���w��0M������v���\��US�B.TD�w)�[�e_�����B��Έ>�*gx���mn�V�8$�q7��\�X9�fj�҇4�E�Z��K6�g�l�
P��@�w&*�\A{n���ϛ.���$�,�����2�-	�Bz���6�'�OzH��}|���+��{h鐮!EZ�����n�CBE�N����.��FDzA:�a��Z�?����ֽw߳��������QXvc�Jk�A��+��a�R1x�0�`����3c�͑�5��[<�͞8=;y>�H�:�`��icw	����ӜiTOwX�<�)s����D�p�#z\�p����O�LB3�
B[�@�N��_u�����qÕ:�lD\���l��������&�����)��X��G�"O�^��7�EUT�2�@�z�7��v����&���u�e�t �¢�i�7J�*��%�M��j�mf{��ppp}�3k�,�w_p�y�į��׍��=�.L92�-����"�I��[����~���`x�Jйp�V�ET��HQB���n�@T���>��]�|�{m���H9����_M#7^����Ui�Zna���Ye�gi#����,&:�qC�dٟf�-|	�Z�2�m'T\ �zD��o�5�þ!�@�A�w�N�#��|�xe`MA���x�Y����X|����aa���kC3�^p�իW{23�Z�!��ұ�IAs Cg���Am�嵪I����@����H�im��^�u8�N{(۳��4wK�4{��s7���i�p6�h����S����ki����H���KLσB��S�W����[���f5���.�~/�c~���ҞS�׏��U�h[T�.+<�ߐ�����|=�E�P#i�Qg����BI�&���2je �ŤĖ���.�~cl1�i���J����잭;|��LE�'�R�&&�~/�<D��{���I��&:�%�D^�r&�E�w��5�4�O��eFjk���Q�3���kI�xc�c�b��ݫH���\U�����h�\�gpN���&�CS�\�R!���i�U��^xch5��|�nZ"�4A?���=�7ͦ����b�:gcG�Y-�&s�㫛A���xo/�܆���$�]Ώ���4ƨ3�#};���yw�Ӥ�ܴ���'a ��5��(��W�Q��Aj��ښ��Y(�nd���-X���dN�äN1E��N�F�~�*G�X��4ۨ�OᏪ�7pW����/�_;���ҧ����L/
�۩_<�ϫ���*��?+�*�-᛭�(8P
�{/]���W�nˣ��T)�䕫�NWћ�M�\g��������ESޗ=K]��C
G{(����?*p��w�ט��7Ʒ���>J�}8*.<(�;����Qצ���`�qu������!&wѻZ���Z��TUNmL_K�N%{W
8���w�h�w�aF�9O{��J=�ǧ��틗/�M^����=�;�ي�	�.3���t��$�҄�H앜M�=��a��.�].���s^�:N)Ǭ*�J�m��C# s~Voα�y�j�5��C��d��n�[�C��ϧ/�_��\W��U�×�X��1�ׅ:I�����%-�E����үp���t�*^���,Q	= �&+H�B��E�=�����[�*�;���x���	����J%�"�����/��~�USO�N����p3�S�A��pzNݍeXT�����z%��ݺ4K��I���zP�s�]14[鼝]�|F�����b��6?��*�D���-<��5����SJ�ɭRã1�M��6�_��M���\�|z��&ъ�f��f\S�zT�� �X�q!>����v�hh�2�
�/G��$�j�u�2��Q�^�{�YG��sM���:������[�Ki�=�~3��Sc��~x5�d�����e�q���M�te��F�"V�Z���i�ܩJ�U��k�⅌�]��= �R^�$hI����ROآݡ�Wm3ƅ�9L-���ض�f�e �Yؓ���=m/۪�wý�״��v�_K$�M'��>�֬��-J�~J�]KyP�ð+��z����c�	���donB���%�;׿#�'^�sԅm����Y?zƒ��`f�vo�3 ���7�k�A0�&o������wAc�$��v񑬚���TɅըK�	�5��RE��	;+h�6�!$c��P���;#a����'��^:&�^J�}{��)]��G� ���w�4HQ����NV%L�7���C������;ߟ�x�vZ8�}�D��������Xr�5���VQ���%�_l���[��,���r����_�Zo�ܮ����7��m�E�l�.��fg��N�!r��vK+)*�~f��9멊ss��_�+�����Ʊd 2������p�+�&wjCM�o��Zή/ó�煽$�U�(�3�#I�T�gU��G��/PX1х�YB���0�|Ԑ���$>B����V��ݏ�oP�=���_ta�߯�ޓ �I�ùx��7u�$�,Ϭ�*xWJ�6�K���6������n���g����
`m�bؖ��?�_�?�)r�a\ƕ��`�1��.��k@�}���NW3c��WM,�}�O��ƭ��bw��y|0,3�>/�d&l����b[F�ֱ[�c#5�c�����a��W~�~B	�k�����B��ʄt'�@aE���g�ot�_"��*N�L^�����Øx�.c&�/z\Yxlֲ�Z�m�@ID�����U�H���ñ�2�9�ʫ�o���)D@����P�5J��{���7���`�D��2�n�����7ƚKH�-a�c|����ۓ��a���/�F;���Mv��}�Bw�*p�}V����=��j#����O	�'�N06u0w�Ș��#ǒ��>�k��X�1B���3w��|���v�첖{)
��9Һ1�^�-�q���x5�I�",�ӄW��a ,66�� b��f�I�t�}`p�x�ޒ���h	�KG�7��ύk,y9��X��Ǜ�_4t��ʧ.�9C$�d�kp� ��\��z����-4w�Ij���N�a��?$)x�{�9�"��)���/<�jl�X1Hҳ�(�+�o�s�Eگ�q>-:ڟyd�b�".n+�EHR�[��ە��S0�ϻ��Lo�u�m���AzXԪ�'-��X6Ϭ��'��̧�|��=4��.-mRV~�k#�ު�s!�7�ˇ�=E{9�"Y���t�G^B߬��v3mu�$�oO+�ѭXt��7l�(��1Ցd.)a0�EjC�/��.��g»���7��ǿ�T:z�k"�$uz/�Z�%:���C�4���Rg�"�FsF�i��j���E�
iq�]�ϸ{��	�P�T1����}�ΎŒ=�'����i�S�*��5�}4��2Ԗm��d�/(QHW�XoA�Q�5aS����-݃��~��3��������s�ɾ��O(³ 'B��"/���\m�y�����&2xN��N��I|1����G�ߎ� %M�J����n�ѷ1��	$�O�K����a�d���+m�C��e��p~!׭V�����h�͚L�b^��(Χ%��'xE3l����EC��'�Y72��%�d{�_$wu�ǉ����M�Q�?v���˙��o3)��1��5a<�snn��hTCE��f4ǖD$�B��aXZ�$���Y�!eT�c`Q�������$V���x	Ur�Z�/.�ÏşM�T����a��0�;�}�G�$�{�����|v��r���t��2�j��f&!���7_/��N�I�զ�c6��Z�шf��br����F�5C�E��w�?��}R�0�����H�Qs��G<MT�F�_�}��N��:n��� {���IטΔU�#����i�yR̕y>�r�O��j͖'A_�
���|��:U������O�L�\�O�$�Ub��kt/�<��7t��|=��S�e�r���Krp7��E����_h�Uy�fy��W"U�d�e��[�פO�4�%�]�cC~\4K�^}�/��(�q�\��ȓc+6�]�T��BX���,�$�aV��U��TM�!�To���2s��Jxxi�xN�>���ؚXp9]��*��U2��Y�/�Xf�����ϒ[W=�`".Z�YQ�$:Vkr��u���e���ՎG�i������n�a�F�mp��\��y��Q*9��h��[|m� ���4��� ����
�,/��?��_�)yH�r2�S�f�ģ��1f���h��fun��X�Is�tة�y$���zS2[
�[����GQ�t��O�����[�6���>�f`\67����0���sqf(��W�����R��׋��W,��+����}s�S�k�Ⱥ/�;�s��t�V�� ^�H�o%��m֗mCmy+�iY���RU6�����d@:�o�}�6Ƕ�d�|>��yA�Te���k%9������%Y9Z�J�����dv.�*u��Y\���q8(�d��������C�k��<����ѫ�d��s=�sΧ-)��)>�L�@�g�A<���YL���h�0wEnӳ@�FWSg�?M���x�ה��~Վ�Ul����҂���HS��RL.��n�1�1n]����x�U��M����rΊO���Ѭ�	��a-Wsw�ok�~���])�L_
�������k�=�4��6�9���
 ��v_G*�z�+ODY�hr�<5m��G/�$:L"
2_�#3
����Őq�Y��v���!޿�8��mU��O�� =�qZ��X`�f�w�"���O��O a]"����N�A�q/&��|�>=n��Q?�=jo��}��= xeD���,�^6���9��֬�&���&f�\s��{�b7`��W�,\u��H4eBy��1��޼N��ΪJj�z�.^ ��^
��ng[ϋ��,�����,J���J�/r���M����R��MkR^m�E���Srw�
`��Lη�Y�+���m"u�� n.��v���?PT�7�G6'��ݫ;#-?��e��'�K|�`p1������ѳ{��F��tMo�Íh�u������$/�c��A�x�@��=����	�ö��=�4pcߥ�Ag�������F=3�b�5�$x����rB(�9ǆ���=Nh{��	Y����$�F��dc�@�D��.��5^+���񷓯����d���$���l0O�0GKPvCB+=���t��|5J�E8Ik�a7ϲ�����2�VI���I}�|V+u��؛����{��+_�\.iN�!sg��<�w�n��^OZxNk~�P�3!|�倈���m�tv��y<�V7�`��ISڴ���S�w"VL��Ve�
�ٝML�5&|���,��D���8�Y��h>Jf<1���Yw�[i��d?�w�ưB�_������KǄ��F�(�X�N���>����{%H�h�s��k׋S�E'�x�E�	�0%L5 �0}ݛ%��9#�o/W~�N�?���=K��<5��{瑵�B?7�ȊOs;3Od�� �`s�͘��s��*)�^ �}f}�MD���uk�H�B���_(��.
ɺ�����9�&If~I,) 5ĳ$��\ ɶ���CǞ!ͯl��NW:�
5O	�9���	������"tڃ]O���{_�"B(c��%�5�޳��h᪲��P��\P�:��8�)�L25dt�H�I�L����}�����9Q��+����֘�����[��^AګGA�C��@�D���2�v{�4�΁	."A���棑��ޱ(�\Mg{��l����b��:ӹ��3�4��S4���02�J�#ɗ��f�Gcs�i��K,���t`l̏t��h���6�����'�$�3�P�k�Sf�B���Nnn��k_w�/��P/%��)� ������ձ�Q��ح&��p��I�)���Q͖8�`�����-[9��}]�?]�?:��7¹z��	�}�M�W*PV����|{��'�5l�sI�\��{v�/�Ӫ᥻��l�ї��d �v4WF�f�	�x��O���?>U����6���[KW�o33���gX�0@���C�	v�VÛ����9�uht�J�gΠ��ⵖyt�{U�o�y�v��_���- H{Zp}���A
���z��w(I`��g�IJp�n�_��U�n��m�vw�/��S �/�I��bI�b��(a�.*���`#�y��B��x������Y��� D��2O���5c�^��_$=w^��b��	'���/o�G�+�����s����ݠ.D���O�+�Ty$�ƥ������R�M*d�8'�����C�[�<�>�R� �#�HO�/c�p��Odrx������zhz׫1Qʭ�,�xq��� Z��Ɵk�(���k^2�k���45��M���tκ�$�O�p�v�<m
x�m��b�#�^!R���T��	A���$��ަ%3;-�א�-_���K��S+�I�w������I3�՘���1wa��ct 0sF��|HX;�&��~�!����m0y�5r�ة/�gO8룢�b�
�%����C�Ӿ}�#����)��5)@X
`6y���V8S(��0A�?��[�>���j��������Sm��M�k	��OY?�2Sd�L?:�Q��dkE����Ü�߲��r�Z�mav.1�-��Zb���f���-��9Y����Ȃ���b��i*G�,�!�)Q �7#ʨHe�R��*��l��9Wba��(�,�ƞ8F<�;q�O�cS&�;Mځ�^M�n��e�K�C^���bFO��O�K�
`H������V�v#&]�J���O~B��p}����YX�[.g w0z˫U�6=�h�»�Dof���p�7��N�<!EF(��a��9�˛��hXGHj\�~�_v��rub�:�����Z�ټ���l�EV?���Y
0p<0�|�}����,���N�J�{桀u�w7 2a���}+?��w1;�d)w�Y�}��I�9��3���,V����r���|}��(-���k'8|�U�ӳ\=���{���n�����2'5:��'��DRQM2�y_��G�i.���mG��ec����W%#�c]J��\���C�e������ݸAч*尢������L��4Ν9�>�7�A�X�ô-�l����e�,fh����,�H)9�����2��k��Ҫ#2ɻ#7���^�S�m�}Z��e�=��Қ��i�s���)�öC�J�5#�{���tRp*�N��!����8C�<�$~Bpcﰋ�������Z̩���+��c�~/�W���#x�@��q�~f��؀�[y�|���s���I:<?��b.�a�g���?'�`�eɆ�gҢ݆���{ t@� �����)��"]�GQ��t��Q �QC���Z 	(��x|�YΜ���`��ѷE��"�(=B��T��3gH����2 iݺē�ΉeC󱋻�.A�%
5[�\�9}�
"wmuo��T��� �U������I��\��U��X=����0G��:��Y*]�-��븑&���2K�����䥴�qr�l�I���?���L� ��6aџ�)~�����Ǡ"Q|��''�C�·:�d-U�h�aC�)t�t6i��FgA�O��<f�RsC���*[����c�K���J��c�Q�x�R�鍠i�B��kA2�3'[��X�q���.f���|���Q6�,KQ�� ����7R.3h�3^xr��u���O.�����ܰ���eH� �*��L�_#`��1��˭��>}dG���<����m�1)4zH�6����`o�_, �������l��t��t13�9=ob�d7������J�ɩ%T�/B7��r�=oձ��mh9s�lKv����뻀w	q_�������$w.��n�_�(dߟ"O�S�n�A�P�j-

�v7@�O�QQ?���E˕����N���BN�욼����
���vf[��V�A����ח�oÚVӲ4饬]���3R�,�q��1��R����;�����TӤ�^��hN����mٮk��\��n�����PƊ�	>cГB=����Bz�%`����NZ�Y<��b����ZZ�QX�yQhl҃Z~f�b{�y*H���)�J8kT�� ]j�V�i��?؄���ŝB H$���V���A	-0.g��_2ƴ����������a��c r�[hTB�&����ma��.��c���х4�]��9;�=) ��k"dEJ�6r��.�!��e88~tl9
:1rHޅP�����}5����m��+�W-�AJ\�xo��j���b�ǩ����{
~��3�e�M;�����O+��\O����ɰ$��]]�nF��݈j��P�%P�h.ʀz�\yܐ|��-)�,���1y{�F��2�I;�]�ˈu���B����P�g�I���ز���p��L��C��G���3�<8N�|��~�S��d|6�ُH�f�f�Bs��V�|��0/���y��+��W�_U�91%[�5]7_6��%F�u�8}`R�hhR�꫟e�� Me!����Y����_1���!?��׮�k2��G�O��b�`�z�����|ɢns}����ZN�m���]RN��rkΏ�Qfeta�v���:`��"�T{3W���s���f�f�2�k�W�%�b���D/)��J�� Ub^�lb� f]hc���e�^-u
�h�JٹV*�x�8���v��e:��ve��9�c����;�e��^9�Qb����I`M6�c�y�����=�+M�ȷrBy�Ο������pL�5]�S*ǋ?����Yk�M{�M;p�����U�@eaL�����\���)� /t/�)ZK�}�~�w&�Z�x��+��Yh���C;T} ��N�
��ލP}�`\��P8�2+d���^�Sԝ1i�=ƾa��T�>�����֘�ţ�X��&#`]I-�>�Z��(jQ����&��,Iw�zn.�-���㋙X�4r�n��G����dd��t���O?��	7��ڙ��$�Pj��o�	P�E�E,�^�h�?_@��|��ߑ�x/	*�hP�䲿W>�oq!lAu��ő��(��x&&O��$ Z?����ඬ���k�͓OgjLS]+����?���f�����\1���B��߇l�e�.�?��Dr~�p�$p��G����k�@а�&s��%y<&f�+Qj�Q7�t -��!������"���Lʆ���P'��2zt�熬���5�3�\a�`.�s�c\��EG�7��OL��p�\�X�T�}�V�עj�FLVA�ǀ�-�"���,��DsQ��q������B�Ƶ���5`�J���8�j��S�VZm��y�т>m�=�1]��ݦ.k�d���[9f5�"/v4���F���td�mQ�i�중� ����KN�ݵ��O4{.��}�������N�.,���>�`1��<�z����2f��F`V�zcmm�<��ښ�k<��/�$��"s�,�wE��kŗ@��	�d�v�5_��1��,��_&ȵ֥*ج|[�A�ZwӐ���"�ߖ�A�9w�S�����s<0^S�{[�Ź�&-��ˠ����ɼ�������Sb~���I���8�Z�s:�Z1\�9	U�\���)�̞���4�A�F-��)���^�`W*}�:�E˧-��TO\��T��F2�����������b��t����Y�5�_a��y��~�
�Д����Y����^tH�;Ĥ���u�0�&��%���B����EW��{��Zj���9q����-h�g�B����V���2�6�ha^L^`��F�Ty}��ļ���
����ž�eL��r�UH���2B`�B�}��_&)?0��k65�9Uf�~�>&1?O�#ָۨ��}Zj*�a{�i�Ic������T��sMI��5�i/)�?��Z��W�7���,���;r�?�g+8c<뀨#���T-�S����5��w��)27��|.3u��S]3�}���z���`�]S��և?���[q�`�:;����C�*���p?��un�B���܋���ŀ���Tqs���"��&�_I���M�g����e��rQ0�!A1����&�H��+�M�}h���f��Փ�4�dJO��G.4���FhI�[�k�9&�������������M*�|�k��M�P��B����nƴ��Oƶ�5�]�~�ǌ>�D����v��i�N@)_��t&iR4�w�+����i����\��2�k���+hlC3�W>r�P�M4�,�eKCj�?S��e3>s�$�����Z�w#6�W\ו�X��,/�u��sg�����Zg~�*��o"�+�e����+Q�$�!�]@�WL1^����%��B6*�n���򮽕�o��$�TE�J�=�C`Ž���e����R�����o���rj�8����n�xL,�>�uk�.&�Ux��[�v��W��9N�Pg�f�����#�9b�՜4�
su/��-�ގU�, R�cX~GI�t�gG��%:�r�]:g6�M�P�%ۧC<B����I��z-�R�C}b�e`Ʃ2Ml�E�O!.J�����������q�����D0�H1�C��Mo\����=þS��'a��z��.��.H���"%�NYa�$T�4� �ٻ%P����~]���O*���B��<r�j�U#�Ez�K��	ן���/��pJ��~�s��������vi?�H~���`ع`�b�>߆ʝ[q�fj� kҨ��|/���:����!J�v������ϲ/�N��Y�2����A׎���]�5�c���2~l`��TY��� ��"�����
��AW���<�ЦW+�5����GN���O{����%�������O�U���ё�!��<gM�����-�Z��T�;��Y2)���"�M8��bg�u<�Y�D�

��!-��:�m+c��A���u��ί^K��9�=7���#��ȸ	�+��Z�U��W%��J5�m��[��t+����~3�I��q*�mǎ����{{�|^hq�JF~}�]�Ujοe�q�UK��L����S�`�2�K�fG�'��������@�k�ݰEuh�@�IV��$ʯ""�-g�����H �n�Q^���ul�E�hS"�� IKw^,�Q���oo�����x�n�e�R���T�ܨ���X3�����Hx���;�HQO��ߴ��<�|���M�M�h�2�S0�:��H ����>c�����R� hqdb</�N�\ʨf�)��.����vh6�f=��S��[����&16]�WR�!M���16n� L�x/�aob�"](�s�M�?�&D�2��Z}����_�R�۪k�!R���[�M_P��	����Q�4V�)I��Q���$M�ЌȆÆ_U�66�&I��J��I���o��z.5Wb�V#�Dj��{����/�y�!��H��t\a���5�r��\Y�e����|���ĸ��;v/� y�$s�K�W��_m����)?��ɖ���`��3�$N�i	���M�Ts|��ނ��v~�=�&Q,G��=��ugY���8֋�]Ia��8�J�3�5�C�dn�ڦ-�;��[�X�h��Q��_e:��ɠ�^�Ww�j1w���[,2�ǽZF��C`>���C��ſ�\j�;7�G�.|�j��_R��rOAu�`�* �"���$�![��,��QUE8MI���FZh�6b�zBB�^�X4�h�k�)��{��r�,w�3�5IO�4j���:]� ��`��+�,��Cm�4�l۹��0��F��ʲM$!�Ы�;��-+u�!b�# ���t ����`n���%�S��b]P�P%���)�C��o#�9E��f�%%q;&��Em��Q�:\?������x��� �=��}J�6���v�ω�l�k��>*lU��^�Xr�Rj>1�iN��a�Z9�?G����y���n䤭�D���@�Y�nϙ�`�<yg8�@�מ����[���4$Q#�t�F/!e�*�
��GM���E�bt;�i�lV苍 ��{s3L��OJ�c&/D�j�Ꙕc����_$/���r���v?��Ҽ%�~��������O��:��E"�-E� ��t�I?v_�����.���a�~�����Z�͏���T�R
�̥֪������x���~ĝ�L�3��AF���77�w��T�z��v)+6n��=]���|ӵ��$��Y����6 ۺ[�hx�xq�r�,�/�+�1�+v��<����p�'?�L�2�|'lVz�s�zjfy�	V�{�eX7b�w����4r٬B�����Z�<�����^z�����<��,o�+�I����hvn��� ��?� 7�p��ڤ�ܒ�Z�0�aUv��V���`���C�G����qM�yq�CD�S*�E(���	�_���s}�ZflF=1�*i��n��h�;D�n��Ɏ�4�`���a���:����s��+��WvOLCBNy3�"_��ʽ{8K�pc@�Q~��D؆����)UXO��;y��|��T�r���Ym�`H_��(�Btx���؉�s4���Oԇ�����l�G�B���p���d1��(?��f1Yo�� ws�r��&�����@�f�g܊감&��oR�����<EO�>4F� ?@������o�i��ݻ\��F��m"�^C�Naq��W]����H({��D�'2����|��/�,	�<ׄ!H�T��.L��d���/1����vH�E���q��Ӹ�:v�y�W�y��D�({t�5�k�%ś��/.A$hq��s|�����F�g�f��8���#��+����B��p�	#���~)�S����_;����6%ս7�.��|���J���%Y����Z_���$3��+d���%������{��9%��h�9��J���t}%�Z�<L�GpMWU��#K�	zЎ'ʢ�zh|aQO�����wBp3�{c�n!ܟ���Ϡ9k���# ��
KrAu�-�R��0�XI����W�o��b��L���ƾ/	<�+�N�I���FYi�u��]S�֩�U��A�.Q� z�TK�9����Qp
)�hߣlOF���sΪg�nG� #�i�A�y_P��%*�
�=퇫��W,?��Ѓ?
^͞�)*�O@ܟ�
VI�k�Zz|�ؐ84w,W�	6�;���<GhF����^�ר�}@��9jС# ��%/�o-�����q���������g��Q���|	ҋ�]�8��)��,��KR!��Z�Vi���Y9��m�� ���	�
h[�[U�c#3<>,h�SΡ�S�x�����v���Y�������=/U�c�,F,�[��8�����~�h���U���e�K�P)���qR�X�ԙW�%�ir�N��ѢFN�ngjs�ˆ�XtC�-)���� *��o-�8�BX�A�z�`��<����2/15��ֻ	�mV�@5C��5O��nB�Fz��o�g�p4_'2	#F��Ƴ�N{� �����a� n(�濊������3�> ���_]a�M��1���\xeD��C2O�m�o���o������ց�&��[�ި�> �I�Ń��̹��ˋ�o�\�HZ�a�"�dޅ�,W�%I�WZv��<_��h#b�+V-�:2K�gË��$
X��n_��f���ȭ�(�񿈉�peg�r��A�Ҷ~<��{��P�ԅ�v0�rb��44
ș���ic�<3R^��çs��:���Q�h��oe�x����f����@�7��ם���YN��s�T����HFuo�8�o� �����9�\ru+�n�?�Fπ���,�}-��|�px��.���PB���\r���w�}*�e�uKTVAw����Q���r	����#�[M�2���楾��G���ߙ�7
��¸��i�4�Ы�	�]���}�oIUq�&�Cxwj�^�����s�0�s{i�'x���
�t�>��(1���4�K5g�k�e� �u�������{
v]u����ٻʧ�ћ|�S�Sn��3��u�xA���柗o=w���z3�ӓ�ďs�s������!��ˆi�iy��!&B��$�6�J����'	H��E%�o�!�"��DI=�>f��c�Kz��r3�`cD���������5��iD�^U2hۍ̐�����*�,'�U��&>Ƨ���:<Dj˲C�H�/�)�U5�QR ʡ� γ��vhj1�\�oЋ��m��F�_a�?ڔ����J�*��^�����[�Ko<��o�2�9V�|z#͗�ێ��J�h혯����t8���7��r�gg4r)���F�l��_zf��w�b�)lO���%
�q��i,B��u�s	U�=&�*��so��ci��շN2mz�#���ixX��֗0����e�A��_�sNOTf��J��	�� �)����=�.=��	xq+_�q��ۀ����U"��Tẁ�
�"�O3"t��B���@�8�_\9���Y}�,Z��j��,�BV'�9!���[��v�s�'���3�Qz����с�z�L�Ag��ܴ�ߖ+�#Zi��2��U�q�X�vh?X�攦�nm�m��ĭ��jkO��wpS��JD	_x56G�'��O�^�h!n4{�Y���ח~Je�|ER��=*ck����F�ѽb��cE�[g�_ {��i��z\z'� J�� U-���[��B��ŶtM�jᵦ�;d�� ey���3��λ��
�F�9�O��1�o���Ji .s�D�$�c����O�m��W��=5�;bR_�h��͒��y�J�H�o�Ф)�����J�:*�^��V^d��w)%8����ٍ�m��V֪[}"Յ���d!����Ӄb�ʹ<�Ww0��$}9i�*]:4h)jf�P�Ի;�����	ky 8��3�A�c�oB�_�{���9���>v%�h��|Ǣb&節Y{�c���YQ��e)&ԍ}���ҸC��UU��w��9�/�2����z򭾔�I;"ɤ y�Ab���/�/Mn������OFM���~�yܫ�"+	���n�R���q��+�غ�BM����<MMxR�/6��+U/���P�wA�#�\����gw >���na�i�F��N�����7�2�o-ɅOK�^t���˳:x(�{�սV�����[�����K�xv�<�����|����L׼�4��l�ډ ��8�6q�=t���is��/�y�ˏ�N�{)���ω����ܙ!fu&2���6����X(b&[�s	�ZT{s�o�0�Q9|�V�?jh>���R�I���LL&��`���g�{���bp�j�8\D�~�ry�Wq=[L�卻\ ��;9Z���JA��d�jL�ж����m�&h���Kpr��yÄG (�7�|.����n�\F�;J���i�k���\�W�?q�{�	y��t������L$Q��JӅ�j��m0���ʩ��A3p��
�"��`��m�`�-ޠ�����t�Y"����v��o�y3��p�k���r:��f���EB�E��F��	g�������ח��	V�z����>g5:������8���C���ڣe12-�.	܏�L��u�h�+���Ϟ:�u�����h�h��@��)3�����)���?�Q�q#;�9��F˿��L^:~�z-�����Z8��&mCڰ���u���B�smn��q+Lņp}b�����<�a��|�s�ҽu˿��������g|X�mi��c��y�"�-��0�PVjn�i���9#w��st�ӹj7� �Pr��L��,z�u)��_�
{]F�{&�$	=Q��2ׅOq�՛}`%!�p� {�����|"����B8g��@���E�1�Z�{$:O�<��٦�r%�h�rIȕ�Yd��'�lne.������6w�R)���e�2��#Hu�Xho��HdۂC}\�
AsE�S�ž�JK��}ZeՁ������.I4�r��K�Q�c�nk]�;42�朳^���kp�~ߤ�M��W��S"rh/[,���Q�w��l>�]wE���COv�8iZk����î6��)D��"�S�d@���HgUo˹�<�Z�2�̪�,�O�LQ�Z��g@$&���=�pztv� �� �X�Dm�B;�Z"�oMk# �|k��x�c�p��	9���m�g���%��D�2���ʨWb-=i#��Tx��_I�M�^D\쇊�Р�ށ���Q����_�q���`|�E*�s�PC��H%@�éDV��}��|ȟ;�P���hn��)��}��LE��N���΁�M���}V����|��鐎AiPJB�!��;�KBA��E:�k�ZJB)iQ�a(I	aPj�^~χ�_x������Ͻ�^{�u��@���M3��iT��e\߯g02�73?z���<�'�pÚb�R�x�SE�9~��\+R)q��ʼ�Đ�RD�*�~0��(k��Ѝ�p�h��{+���y�ۻz�mN��s@�b��x�ރ{����C��NB�4rY��c��0uAqm%E�F�=�:4�,���ݾĖ��O�*I�����_�e1�.H�]����?`�M�\�jx��u�'�	:GNMV��<<����ʩ�D@k���[{��&Qc�#=U3=o�����ηR]ݔ[ \�_�}���L�<�~�O{sts��
3޿�Q���� � ���~�蟑J[x\�=�]<���u��7z_�c�L!��F���i�W�F�#���X�z6<���R	�@�T�ތ��4�{PK7FU��gM���/���\r��yv�Y�8#��v�X��!���j_M�4ŭ��N`Yh�����gW���J,���qV8%�>vЂof�e��5���ζ{Z�3v ��>�yy��*�k�&�����q��GX��fu�g��A���������d����.��c��� >�?4�������:�Qb$�X��k��c�Q�qϛ�H������f.��`����?r��=�3\����רՐ%֝KX�]h��k1���k����:ǲ�b��3�����Z8�a#t��� ���Q_,B�ԫ��Xn��j��i`e>55��*���{�.�:����R"L�9p�ҝ����S�o
.���i)�S�I��l��!v2g����}n?�o�{�T5�P�לU���#?�IOHݙ��Ev�ߪ�k����x���`6�����7ь�hY��$[D���S0�E_�&k I�.{>��"��ӫ=J.1��e��u�ۑ��\wJ�uq��P}�&X��=�>�F.�]�h�5JD̄W�-���cxt�P�k�|�����F�e)�	n**�Z�D)Ir#�[cKz�ځZY6��9�4
���8��n:�@��&Ιr��/7_�d1�ʤ�(B��j�):ܳu���s�]yp��J�%�oFϨd�3r�u��m�(�Ҁ��e�(���$��y��wB9�L��|�5Ƹv����aAE�9Z,��z�xf�3�?�S_
�.�� ؐ�[k��Ĉ�Ļ_Z\|IpP^R���yT�9h��ʅ\��{��\�_}�c2�h�)���Lyu�&�V��[�1�����[<_�|��]-�5*/��]L�Z�K��i0��R�g���{��}����;���h ΐTU�Yꕇ����Ț��o&���	�k��-0*�Sӵ�LTV��(��?���{�w'<櫫T����?��>���j�Z�2_y�����5����L!�Ժn.g�[�Ig���;mm�Վ��ءr���- <�&�Ly�Ɠ�ٙ��!� �Bi/�6�z�,<.���i�o�]��IA�5I~0v��C�;E�� #G�)S�)�կ�1gu�빥B}Oo�@�������]����"��������s�N��|��z����(�<�;��h{n2{�n��_zD�q�֚�A����Sߗ��+�����g��I7���7��|t�&�����`��Q}�C��K��+�^�e��fi%��%�-2�4ja�����VN���;ޢ��UL�ḍM�19��U�(ML�]ȁ�}/�1�N�^O��}����~�`a�b$�Y�u�Dv���R��M5yq�r�CI�ѤAi��_M�3#�Ι�W�� <�D����/M<��u\��u�իi���5��ܠ��"���)�M�N��1M�g.0�2�ܮn��Oݨ�7�|Vg�֛s�l�=�lY��	�<~���/ޭ##��B1�5ǰb^�)�
d�	},k�N���� ~S�ho���t���K#EE�F��9M�\؋y�M��h,��Tygm+	Bۃw��C�iti?��^C��:����{��K�f��+�,�����?�}}x��Q�3!�έ|h�yN{i>.�z��Ԁ�BR��/@���H]�U��N���\1W�m�me#OD�r�����+Z��q~�Y`  ��f:k�Uɏ���fB<tb��<At!�_mӯ�C���K:���*�e�<��觅0h]��ڇ�=mE?��V2���~Jp������z�V��� ݖ.OKB�}~�!�ms��}��O}f��c��V�C/͔��*,
Z�+�rs��p"��+%������^�����H������,ъ��o�C�7�O�IM�����Yv�37�����gy�q�*)�U���}��{x��C��"���V�zmEz�=��j�m�U�-�/�Ȇ�:	�ͪ��K���T%'&���r�'0�^��Ȗ`��O�����Ĺ�G����x�U&<}n���\'�bYy�����6�T��ʟ5��t"L�n�l��G�dG.��Գ���>�kl�&��5�<�mY R  �ȝ�T�S�?���rh���6����t�|b~��?����N�5w�t66C��G�u�Pע�_��&��	�$7��I��Ƙ���[����L��7՞z1�DW6*X�s��Ǌ'@0�9��@+�BG�u+ᅼ�5屌P�c'#��cX��\^�NR��Xy?�d�j�y"chV�!����;-@���IWVgD���H�Ɂ��Ba"zU����M���e�����I��9�3�f��-�i�25������r����}���;6��d�-���_��Oҙ,t���J���S�U�A��G�z�)G9��=�+�!��!]nf��Zi��N�5�]9�F�d����{r���,uU{��L(��lŧ�%D|�T�Y�\�d�\�j�Af������q6Kh��7>`�ܷ�q�V+�$S�'�{[/�I_Pi����Tdं��p� f �8�L�7��i�\M�&��&PH�hJD�}�T�G��E��.�8m�2}�c���z�}�7e�} �~2�5Uv����YvE��Bc��p��?a�5CN���?}�𔪁�YS�ǟ��:���=\���n��x�5_�1?{�V�׾�l������ܠ^�x�:�Ѭ_b�_[��壽Z�Jb�KJ}Ъ?�ne�­���x�q6b�7��g2��$�sj�%C�E����4�܃��1Ӱ��'���K�d�e�Z[�'9�|�	*�4�
p��"-֪�*q�%�H���V�����.�R��Kd�&;5�7���ж@W��U9����W>7�W� ���ٺS7�)�	%�#b²��U�|�&SI+ޓ<a��{3����x��W��b���p�N�-~�J�9A�:/�_?;8J�aQ���J!��o��n��/,��+�t�{���X�������pXv�95m4 %���r��}sJM��G@+���[!���v�����<��N�V�T8�w�~p��7j�u�e�PQ�4MB�د�����9�3{�WbO�'TY���C�@MC��T� Y�XB0�`XԵc���8*LsW��M�i��Fo���EW�����-�Li�Z��=#w��c�"r�P��EÊ�۱���׋�w���9!��)r�P?G`�G;�nyC,L�#�����n�-�7E��FO��rLN�P��c�j%j�3�-|((�r\�`����C-]���L_�iCN�9�럻�~#��H���jj����yq��U��1�4E�Ѝi�fY1��.������NB&�Lb���]]@x�\�=����{��Ȇۛ�����m]�����؞G�c\�Z���n�n���AG����q�̮̾@���������dM�q�C����(��(��(m?��v��<����A�w[�'��wt��ܝL30��1������,Ʊ2�8��5�"{�`'��G��_�0�,o{���r�ʝ��4�Z>�P�+���J�h#H�%.2尵��`�H&�P���1cL?�m=��ˏ��++9"��q��y���e܀>��$y7�Y^�B�~"L��� D�V��q��2cH�	�E�|1Wן��(<����G������nnr!���7���8��3����B=.�M$��g���tb�r��r
�3��Ҳ?��'&n]o���Rt��d�ͯ�"#�J��g"�	B��hV�ű0qBubӚ�.��hꜧ!E
ם�_o^�J�O9�Z�O���#�y�p�a��h�@��j�W5�rBҗ!����F���;(��փ��a>{0��[Y��*�Ά�3�%����#?5�Ǳ���g>��������j_�%rvV[~@S~J�i�N0����~L��w>Vd<��)zb�N5
���ɶ0�����2�$|��� ��������Խ���G�o���w��sH���v��t����v����h���`����b�_��q$��{d�:���m��s
���q��Ba=�M���^K��Xf�����BtG;�kM���>��_!��n~F�I��������240d1����Fc�/LH�U`�;^gu��� ZLu�����lT"�}�gV*a���3��y�p��>�`�ϠEU�o�G�Y7k,	i�)�3�B��c��|σ(���� zmd�&)����a8�T�l���S�����~��JA��]܄�|"\Du�De?���n�t�M�@�Sg_�7`��AJ�K��[�1�eމ<��а�����R����9@�ʍ�5�/�d Y>�u2���'?�T]�wn�Z> B�c��5�xfQ�8!�X���N�|z�qG�y8O��w��Ψ�>k6j�,40����=��|Pn�&8���h�:0A:�SQ�JG]f��JE��p�O7�D�?x��=�a�^��e��Vo���Rߕ��ո p.�n�_���d�0��)��0�P��cz?�l�ߗd8FIM��f�g���q֤�Y���{j)k�y��Ea�I����r�����]�h`[z^�e�H�=�J=��w��h,�V�z����DR��o�����n��z>kec��iJ���X�����:<>v��qh��t�Q��#��#�ټ>�ޞ�s㋳:��g�j��iH�]�fqu����=BO�qKW����ϟ��V��JL(Vi���qŏI����:tӤ��#�,�ūeY��A����x'����֩E9m_�gy��z*�0���k]_Uq���>hg�-+l��LnҐM�A�����D��ZO�S���5�[b
�;���{�*���^�n=���;�a:ۅƴ�(c�~��5{�׵�����$p}Ϩ�@z��7�'��=%_W�$�κ9@���J���UH��Z_#w�����r֖��$����`���/ݧ��z��BN�]�(,�l~1�lD������r�������YL�F?�T?3�Q�Mdn�'_2�)�\�6Z�e��R���L�6�Q^���x��aG������YeY(Y�(t^���3,�8��N�nVSK�=���֬=Hg��]��<���;�?o1��칀Y�������\��Ud�� �!�����9�� yb��LC5i��b����ey(��J~��2;&-4�Q�%H���W���N�~k���[��'{u#�����ʒV�Oz�ޏ�A�/���^~SGx.F=H:��5/γ���P*}Y�a"�ml����a���m�T 1��6Q��7w�������<�:.;� h�/����6y+����a��<3X�m������#�s)�2��U�'��ǳ�tB��F\�h�����\��5\���m��}b�����|kM�5��A]T�|���<3�1�㷠�6�	���Y�K� O��F����,MFO���Ч��+���ykJ�fLV9��Pw`
���'��c[�%�4�Y��o��_t*�U��  �l`iW9�G��0S�9oY��Y �?>v.��Ɯ4��t�;g�6��+34D�.�m�V>� �5s�/��׿s-�'���������Έ8�w�����|��\���#�`ɿ@����l�E��<'w$-k�ڠs��;�,���4�C;[M:�Br<u�ۙcM��Ҍx�B8*ʄ�ʇE���d<�tvҵ�cЇ(0럾�؜=�G�"�B���ݺA���.x��S�����f^��I� �U��77�~%��&�Ve�J��^p�^��W�,��k_1drn�\�*\6��+yM�^Bb��*z�q���Y�l��؎I����hw�kǓPU �%[Uk7M����?X�E�\A�'��_v��Z337
�c��\�L�/�Ɍ��J^w$��e}���L:Б:��?{����_	<�FXF�|i����z;����tI�7���Z�F�N:gȿ�,۾�(��� ��t�����O�7|��G,�}���W0i�Ψ�Y�(&��9�6�Ĺ�9�r�Q�>�P+X��SkK�o��K���O���턅T<�����[���Y���1s��E�A7^T���RJ>�}�P��>U��阈0�H�S-`4bǢP(U�ޒ�d��N|v��+<�Zf�f�zsr��ٿ3q󩥌�
X�+��˩~�/Y�����!�iSX68�)��Q���RI�1���Ȥ�|��?�w�bI�ef��)vP� v �k���9���X�B��{Lܧ�)'H��%3��XRD�����#2�U��g��o9ݵT��8�Y[U�^!��|�+%{�w߇�T�Ve�@p�<�T���y�(K�G��Ɔy�!�����ͫ�W��$�� ������Y�	5_��9���%�o�w�d��
���M֨��_� ��8�7����4]be�v`���I�:wu��^EM�������U���{��X��� ^xţ��0�p��3���꒯��O�R^f��s���(�V
:�Fw������ٍ�
�ũD0g=�IG�HYù���jm���Y�Z@���.�l���Pn�~��ۗ�Q�p
����C��qZC��k�Q���4@$��U|�s���l�VE��&o��Ya��b���Z�y�ꨮq!�X���Ob��I�@� ��ՙ��A�;���~w�����v�T UK�\ϡ��ʊn����1܉��a�J��c�!���9q����ԏ�P� c�A���l���z�����/�bw)�U�c[��VW��L�!C�3��\�6b��ĶǦΨ�D����Sx�����k��t�s��gg{Ջ�\vv�j��"*�4k���x�,4)P��f!KD��>�_�6���>�V� ��q�u�uyW���<ؙ{�Jc����R�ۮͥ�ayݲW��Ԅe*��8��r�(��g���T�+d5Kqh�B;"H�jb��n�8_��W����+�\@�D�(6�������F�cU)�����;VVW�ٛj�>bv(Ҏ=3�:���"SO\v4j����o�qo-�UJ�ȳf���QH�>s��=�K��f!�l7�5��Rw ��~8�w
#�+�����SӞ0<���7���_P��$���I=k�q��uO���F~*���ռ34_����Ǝ@����s㡴n��B?���*լ��_���޽�7AJ\h��4y��s���;bĞpw��\O�{s?v�L�������LW��� ����B�x����ҹ�D�y�$'.��MC�,�f����x$��t�J]V�p���r�
ȗ��]ReD��Fɿ5��'i�$]��f�O��w7jxYJ��A�͛��do������H�&��/W=�x%$0��4��N-w
,�S{���j�CkL�Y���jA.��ժU�U"�)S���$|�rK��?i��S�u�8��j
PTU�%U�q��.\7����9�����EJ4��Lh+����4f�+���Th_ƽrP8���|�_�G?o��e�u�im�]m������_=�:��QT�L���3}Y+��ӻ0�B>�V�����9��-,M�|g��RS�<FE�Q·{��(��3Q�o���ZQ߿J#��������,�{����+_��p�ͻɓ"Ԇ���p� �l8| ���A�#1�k��w�x���^�����c�x=D�`�έ�K~L)�MLR���j,��QS�ج<�L�'��,sz��?�3���~���S ut�uw��������_�t�99�yP۾f�oz�]��k�~���*˽�-���i�g����l����,w��}�^�o�����C��%	����]�Ԋ4w�8���5�A�r��x^�����"v�����ip�&x[yҖ$����YQ_E+�|�2�_wߝ&��*m�oj6y��m�~ܠ�}κ/Ȗ/͘ п	�?��x�زx�,�@͍��~���g�n�XvAJ~�����(�������oA�k��s���h��}l�:�A�wW��6n�F	b�U�����?j�rV�B�N��:��oņ�0���9ݸ^� � ,Յ�o��]���/��١��B����ʣE��ǀ(g.v��'�8�rO��a��p�W�׉���5��C���� RL�z�_�pg��6�Y)�Xܷ62�ڨu�I�3�]�~��uȷ�{@�ʣs�99S+�mV�� �nC2Ɉç�,���$��W�,b���j����_Q���PHgu������-�W��P7�=��yό���	D�����Mr�KC���E��}�i�LHq���H)~V�b{E@���ff)�ͣBD���cB��fiOFԖ�����ײ�"#��H4x�U9A���	���|z�ܞ���;D�q��E����-���j��I>h����DQr�Ajml7w�ly��U�&y��x��%3�U	�<�)S+)�"/�r
g��0�,HN�N3Oc�%V�Osr�,l�R5��"�t�5�����]˘2o�5v!"����^=���6�7�S4���z)A�3�A���fb�/l��w��^�vv��DT�)�\-��5j��!'b��c�n���S��f���x/3�O2Y�z��{�!��R�'���n�E�8���~��3@&��F����XQ�P� w����*��|���:_�ϩ�ݼTn�� ����5��d8�U�����W߭�152?1��bp�sm���g�'���\�8�k�n	uk<`�����?�9�r����V�e�eQ.he��H=CP�N�luL]��|�*Do�KՐ��㡀�$�=��z����Ar�\�<�*�c$�Y��xs-��x�������[L/_Xx}�
}��]*��iS�$Ł�1���~�KV2�����VVoȬ����%��:�E2[��X=�O����2j��+�!m۽u�f��/~�	�n{r��X5BR�,>)Qss�o~ل��҉�SRR�764|�@M[�~ҳ������]OR~$�Lz�ha��/��:�@��HT��R�E��Wbn�AbI�\$ �� r��@�CY�*�T�^<�	�ǹ���/`lo�����[��@M{��C��aBK/����E������"Nuv�B}���Y&���V@5��vuu�m	o���:�4s��7��i�B�q���Y_MI�x����EV��6��ݤ�m��*,���h&L],jۿ��'$��t Dטj �n㗡@����*�Y85�G�� �����梻k���H�㟵\��$U�=�pn����N/t�Z������g.�	��^~�7<v�Ƿ�G���L)���U1���"_������O*k�k�f���%��C##�j��Zdy�s��d�ys����_���i�e��������{8`g����\�`��J[Ki61Ѕ��	8*9�������a�R�  ���������&�W� 2�H���m���:ӟ��������J��Ϩ�˭���!}T��{�&��ˮ�I����������k�#�bӛ!e��{B���Ե� �˲2}PF�
	�ڨ��5Mb�
k���i��E0�&3� �g��!�2��� ��ˏ���R%����u1����w����r!,7��F�Ty0�}��Lm�9JQr��g@J��b��{����4�����Ί��Uu<��- ���\c��C�N��9�S:m�h�C黇[Z�y��ҹ��k>��W����8TdmǨG�Fj����Ȝ
�����S���"^Vz oH,=]AU�������Q=���͟V�8w���Qg˴������D@r�@$�`9��E�7OpcK[�S*��}u�+��+nƖ��-I�����'\�E��0�R������N��L���V�����wJF�+s��dDp��vL���w�jᜰ��)��Z)���k���P��#����'������%گ{\���O;2��3�qJ8��S���~ ѯ�]����6�.�]��5���9@��7��8���.sVC���|�ʓ�|Wⷀ����]�r����~�Va9���m���P��P�?}c�&�F��V����L��@��e��Y��#dp�(}{���2���X{��3�G�6,"�ǓK}{W|g�S�Ad@���h\s���W�5f����{�}�*U��S��|Z��m*�����6��q�Bt���٬���pԝ�C�л�4�#v�.�ϡ��ja'�T3��b��T��IRP�����i=HG�=P��َSư�#C4W��d:�.-d�����V��FX�{+���p�Z<��H�������A��$3���S��+Zߒ���C=PhT
JʁJA?��=V����f���Ox�`X�ʧ$��
��*��tX��4���ga�%�6���B�L�OW �JL�E�v�zn�΢��<V��~T�hO ���u��P��[���0DF�F}T�-��h������fn������.�!�X�m������-M&տ$����m-YZR�5OAF�4���%\�s]=^�*s m��K�a�^>��#0�������L���4}x������v���C2S� ܟH������%�k>�\FN�ֿL*��i�PAgǚM:���,��`�?�6'�n?5_�R��\�
-� ���%����d�¿�2[Z�K�a��ĩ��/1�qS~���2C���96��\˨��L"��#�!{ך�#�V�e%���LmQ�;������`�2 �L>6E��'��Ͼ�-�����R�
��^��M�_<�"{���������7!�o�:h�!���| ���|�"Z�9��i�i�&��Bd@�׵����̕���N�e�}h��V.����v�y�H�*V������y�!Y�rїsA%s��5��M,���h�$�2ȒIu�3�|OMXFE\.! z�QLk��YL�����m���"�l�d��F/ņ���R?ַn������M���d��E���?�_���K�ݝo��}?�~�Y�1�\�%g�@�9m�!��}�|=�X7��{N'��@D��&s,�Y�׾����n������v��k�8����6�3j�u�
j�t���5�����P;��b�4�Y�<j��5$�/���7֘�0��:��9�����i��sK=�g�2��wɻ}�۵퓮�~%��M"$�v����^�_�`J���E,
o��)����2(3���<��x��(��+�Z	w��&��F����ӿ���DhT[��[���;H7{��P�w3t�/�ԠXb����F>#���d�n>,��𣥵9�Za������*�r�}��i��Kl�-�&Ue=5yS�3��נ�ٗ�RL�Qb5��{ޑ~��3�@�4Žf�=Tgb��;�=̝8��g��T��������1{���S��x�����TU���ջX=�M=���`��@�����J�j�n��v�l5�53w��������W��E>ɬ"�S"�$�N\����n�g%���D2�^��%yU��q�/:\a�~P�A����ǭ�y�=T��3�kG�w���Q1V�R��"�x�\eUS��;���=_��oԉ��a'+��0�ۻ��Z+^����q���oF�yB�*?J5��VԔ�2T���%p�	6}e�4-���o�2����uN��T%��Z5��?gi�>yD��I"^m�hP���&p/T�l7M�`D鋻�����=�}����v
����Q����؈?,����~}���ap��-!��T��(�}�y�[�#��Tt��\�2;V$����v����P�2���]����0� ?���G�6�4��o��u��)��-MÖ6ǲ�%/3?��T*���S��<�9�T6m�<d' �|G�(�c�i�~Fg�\ͧ P���:��C��L�5uS��4lPݗ��+�u+��� �C����i9ʮ��iq
�%&t��r�(�������B�����C^jμRWsJ�6t����3F�[N�|�GQh>�e>K��ц���/�Eδavr�Z��Z�3��$^&�&4�h,&{ h�y��'���N'�i)[�~���9ro;�⬿� .��� �{���+�*M��H������g�dƎ'��Y7А~��9w�F]�VZY݀�`,\Y��S`[�Rt0�tT߾��E��'�����-���:�~�M�y��\� k���k+z6<�li\|���L1}�M�ӥM�e (-)qS�&�?s�z�V� 薥�j$�k��E.��p��{�MRv*O��G�����-y�<�Qŏ_��P5�a|w����L�e��އ�G�Ԓ�C��]�D�CBE�c��=4X����pv�	�*	��n\	އ<�i��/._^�1���Dԉ�<=ˮ��_mT��?a+6N��G&j����r��c�L�̲��\�:��6�N���#'�����:��,�ܮ�4��<F��ز]O �4�VC��5J���A�}��z�j�l@��/$y:m�+h���Q�ɮ�Ή����A�`�_��'s��[�Q��!���Ŭ�	�բ��e		�]L9cA�O���r����;rr�攉���خٿ�${()��A��M��V�5:8%���+����d��G���UHZJ!����))�Z�ڛ���{]�D⧴�x/%^|OdR���_�b��jX�F��?m�>���Xs��8]9�)i�x��ײl�^/��Pʾ�5ݢb�x�;H]~'�_�����x�866^j�7Q���)��=�*�oaҪV��Q��M�/~�x`����;��I@|�D�,!��
�n�Y�܃���:�'Ǭ	���OqO��s@�<��	,��,���↖� x`�|�(�nJ���3�_g�al�}���`T��r-�5#��@,���0_-�a 4�L���5��X0�7���O��[�1xo��ȋ0⛵�<���So���ZB��������� ����,�e���r&7�b��s��<�e ����`������ޖ�w�v�����U!{��н�r��n���#ɍ�h�{�̎��/��;�&1���dM-G@L����+�9��zFq��mkr��d6���?���jϊ��BQ�ab|�ǧw��G�~d���xE����;X�	2(q��.y�ǻ���J��@�&�ʣ�g�h+u�Pl�n5��*�c��V���f�V��*m�i�����.~��`>���$�Qȷ�j헓�f��ID?��G�~�]���OC�l�r����E
�1�XK�Hw���t��WX�;�Pq���*)f������ϯ���M��{���L�����b�<����(lr��G|�$�4T�Q9���9ޭ�g��T�>9�M��}| �Ha�-��ܬLu�ׇ�ބ:�Ґ���՟Y�)�{��,���v�ȓl�+s zjq�hnR�e�衫U�Ǿt���M���on�-���_�gԥT]�e-���3�r�!�:VQDY![����xg��5�E
�;�}�-��7��t� ��ڕ@n� �G�-�������޵!_oQ񲭩��G��?~�Óe�_�}�K��vJ���p��v���5x�	�2I�������M����X�dDq��������I��L�P���2\x� �@�[�L�.\+!.Ug�*���'()��f���?H�Tz��'�E�X�����3ނ����B.�;9��=ad����P���N�{ua���wnu�~�v#�|§q���z¹�����NS�
��� �u#`�ɀ���-G���j�6�Sg�����Jo�⧬��3��:����t!���Vc��a��FaR�~)���7$��{��,wn.�$Ș����O��Ɇ����A>q�y���?ˌ9o�F�O0Y�o�ƕT��e��8"$ t�x\����#O��L�/�a�SCwPZ��ңȘ��S�/��jzU{ۚito#��_�!k�gl��c���h��߸��c���(4�٘� k��WN�G����!�0cf��\�/��1c�s��
��ۍ��[�-'e�z�B?1x?,��zf+���B�1Tƴ�,�� =8�#Z��Xg��`�n��V.&)<\w���@�al�UBZ�4���/䈵�@bd���oy��t{�,6rU���bOƴ��� Yǯ�N0{"&Y�w$ 呿[��{�;N��w{���`�-�\���f�\���,7>�>��U��J'���LM!r��f���Tߛ�~d�jJ�O�	'��~ao]�j�w�87��Cfq�^�A|�/�%�UA�f^��[���
VFc�-�@�^�y�?��Ƕ�K����㔿
3!����Mb+�vn`]!۞�x�=�^��?:Y�~9M���耀�"X��׎>d{���>�ĺ � ��G��s~���MO��C��O��ۀ���#d�����7��5�Y�D�����`��D����Ω;�D������1�,gήm�_�����A����Y��;�dڼ:	���)DR��ԙ�PAnOBz=�I�	
a+(5�^	���65vJ%+�\[��)2O�D���T��##5g�R����Ӽ�y|����/�ǒh����0A�9���՟##^��>F�����#�I�1��;{ۖ�`O���z��= h�@�9�+^�]i��+��0��(��z�G\>,�������9?(�/��������?9� �^lҍsg��0�Qc���ӑ� BwYp?���Ҝb�	��m�����Y�p:X����.~>��5�٪���4N
z�dy��D_�,Q��oG�d䔃�k��
�h���`cÙ�'��	�]\�u㢔cOΚDh�)#H�25�\^p����\Y��\��8� �$+�u����C�G�阳���Q�\���|��Mir~g��0�+;����1!��D0���;�|m,�!8k�Q���K�����/���+�����j��r�g��km�I��oR��|�(�95�0�<���/��7G�E �T��^N�"0�ܺ����(?3u��mp�i5sS��R��n�_3����hĴ�}5oU�+(p9�~�\�l��cf}�P�=G�� �[O}�Z�Iajr���w��S��}�4r
C�6s�'U p�AHl��5;��|z�N�l�q�3�����������ut��֗�5���Ԥ!�y��c���K�
K�'�X&��F�K�g�Ԃ�D��_5�*���NS##L<����]�Lr��vaD&��u�zVo��<V��j�vqio����D�S�yܰ|��`�'~y?E`,��s��afi!�z���W����ɆWwnJш��L��Bҽ��9Faą�^���ueeW�y�&�U���m�9�����kX���W�����և#��D��Yh1�W�n���e��{=L�3Y8�����q�z�\7)�@�ȯ�/W~��A���@w��j��A�#�݌��K!��5�ِ�$-��Tҏ�jt|����mc �9�!�����L\����>��5c.@�݀d��MX��^u�����,D��_#0�&t���O	� K�i|�֓	B{����(/�ٛWT��������j�X��!��ǐ_���m7x�T�O�	l*:K�Ɨn���o�^�k�������P�pU���,�gY�Ĳ�A-�"#�N�_��D?H�9D*B���'k�����,_/ylkX��A�g;�w��2�.uɆf�d�	�J�J��Qɢ�=�זyjU�����'�b�"$�h�n:F@夙 ��+�	�?�{���_�nZ ��xF=�AY��"��"�NWHu�h�fc@p�8�����Ui��z�ڱ%�w�:��Y\��g�Ŧ�|[��?�4��;{S����[���eU�o����(� ��2��rBr|_�^[;��m�\�?.��5���i��/>p�q?����r�S[�4�ͷΌΔ�}�sO�s���9?�W0���NWQ������l�enSY8��E�kC%�N��a/�
O]��	T/���B��j�5���l����꿨�h;��%Hw+�CH��]R��CHJ��04��]�J7C(- 0ė�`x�����o�~>7>�s��k��:¿�ħ<�w�F���'C��ݘ���T���}��1*7Uw�Q�ٓf�u��n���z���y�h���W�ܟ���!�M�?�����D���t�k��'wy]�4���im��Ŕ�"�ć�U�~5R=�5|`������hI��FcDD�L0���{��������R��dZ����1^?��vS�unS�(ם��������5.�,��y���h�{�o23�Dt&I��&��w��g�Ld�s��#I~^Q�>���Vp}�C��겕 G<�e����rs�wb�+�T���f�n8��O�p�G��	�d�������7~�u��N!zt~E�M���{?(�MYTF�O��)��I�F�U&)9{��h6}yC��4�t���L$��!����W��]�e�|�Q��EU�w�7�$(����t*����`��f<��5-�|nۘfr9m鞡�~������e�[�N��i��C�R����S�o'��sl@�d��+�`Ķ~SŜ��א�Ǉ�s�,Tơ$�Au��_�5+0�f3u�
��
�$�q<�Х[+(����i�વ<��c�XD�%}�-L�d�h��eIğ�_�ɓ�܉a�\`��`p�w��]d����3��o/�9��Z�kE�����쁀�I��ߏ?��"�I/��'QВ�Ӷ{��ζ,�#@���h3,���pѣ�F޳#*W,��$D=yXT����^�!;�K�����=�At������'�H�)Rf���r�j̇gǙ��/��Ep:�_�k�w������q�;V��♘�W��b?8�e����{��K�oll]d�o���Ru&�h��+k%/AD�������߃�t-!(��Ѡ�~��w��# �@jىg1��R���<6�]�7b�u&��HL��?ɔ�&6�_o;U��_¤ʤLd�F�\�c٩��.kI��N � }eo�F��Mjh����O���������7G�j@�����$r.�`t�Uo{�� ��0]�T����%�K�@{ek���?_��/k��.��4O�ߍ�1q~�}*\V������j�X	��a�[�L��Ȟr�>����=,�]tX���X�_`��Q�i;�ڑ�$:l�ʓ��ή��7�����\}�4)�'������B�|]��5X���8���܉�M�P�S�d]3W*x4��_�I��� ��@Y��o����o�`��^�2>M/pF|��T��i{�T�D�#ʵ�� |�Eo�L�?֩�ZdX�~���Pct\��[T��0���B�;�$�.��d~唺��ƶ-"j���B�9.���?�g�>^-��ԝhÊ!��L��@�����=��_�$k�����H�μ{�{(݇A<��Ok�!q���4�I��'&˦�B��#�]˨!MK�=V�gFH����T,�H:ݽ{�P���[�A�j�ܨ��	�l8t2o�@�pdN�nI8�st	q�%{�z�?sd����\�u��gg!w<Q7�2
6ggI�p����.^�2�a��A���兿}�Kf~iJ��Rc�P*ٿ�[�2W�c�O~B�Le,w�,n�J/��T���1���`�쉬 ]dX4�z�ʽQ�DY��G�"��Q�)�ư�a|D;�-��2�yc����#�aȷa�ι�<��� �+�$�Ě��y��^3Xj�#���l��j��K��w���;� o-��<��K�Mc����6 �vEқ��f00
��,P�-���c�����������QK��},?s�)|&�~�|~��\o��9�we!�G}}���|ͤ��FQ��&�t�����k�%T'r"�|B{��zO�w&!�����Z��b���x\�|�z�e�euK^]��k���G������xɾl͍0}��l��N����tRk�_����4�����?v�i��^,�x��
��#�TdM՞�S#s�ir�w����&���Mq{\H.B���	� 5M��{9���6�-*	��ҙ�Ji�@3Y�wI����Ԇ�w�!�=�R����6��sQ#������T����(DQ.���ߡ+y=A1D;h�:�u�?�8%Αk2�`ʏ���*^4�	5�]����m��R/7�RlT�,�NH���]����/]�."�Ep=���"��=�:��Pԃ���([��3g�*'S�*��5�w 1�+RO�k]���j��ޮqQ쌐�bF0J��%N�=�?���r��x2
���-��BD�)��P��p��;�䀖��9_*c���U*b-'�V�#f��z�ͧb`"X�����I�Ý����9&G���������Ke����k���0G��<4� p��́��Ka�Jb3/�e�i����;�ue���� ��ٜi�K��BQ&[��ӂ�� 4��mq��r��Y]��O�*�?	2�l���ٌ�YW��r�y�	���`Ȏ#���TT��ڪU�Ȁ�J��5$�ٍ1+;�b�Ff����>U��1
b��K'|��7V��K��E���!�5�4N�|��̈Ë�9m�����"u�ȶ��������J����, ���V{��ő�L/��oLn�%�L�e5)�x��C<n�� �=9�m�Þ��-�	G:+���n����;"�2�2Q}M�'�ʯ�23\[h/x%(����u�%u�yo[�u���ݐC��/�.�娕����"����5����|%���x���a� �
���l�\����z�������
�
)�8�dB1��v�l"b/�Q���r����d����lְ}؈*��j��C3��D��sT��K[��^��&��Mh��ْ����ů��h]h(b�X3��8�~�b�	�A����VB���t�>��,O���%p�|��Cm�z�	�~�%�9��Ћ�G@����H-���9�Qj'IIգ�Go�yX���;�)*���}�J"|�M�416�[�����u�A(N'<�(�x���;W��!zx�7%?-J/�ŵ�6N��h�T_�,!L���$��V~�}��+�sH������w�γt�/���+z'�%����5\�,�Yv���¸��;�R�C�mC?e����K�D���R�Mb� ���'���-'sx=!@;�̴cRTel3R�3BO��#�0P�ȗ�ҹ�N��M&|�=�:w+� ���x���%?[���������5d�f��ũvfV
��Ň�.'|��u�A����<>$��}�)`��b�+�Kԝ6�/��l����u�*zSDy
\� ��A��	���)��Y�LSI�@����ƿ
zי�~1���4��r}��J��ގ��Z�Ά�Ml��a:*z:���G@�W�:Sn�*�Q/칯�VjJHNYZ/�����܆�ߛ��8��l>�A��!4��z�^e�\ې����*hΝ��+Jze�2���v��j[��:�v4�K�րcwa�T���L��^�O��F[���úv�'ﾁuU[��2�=�S��թ��:�_O�+������Ӽ5S��
�֌m���5Y�~�5�������5�Kc\�+�����ܙ�+;P���ٴ���z���j�����lR�>�+�eː2y"$ů�裳��d����!#ܕ �hp1CjC�#��6t����9_N���<ew)M��B�J�rb���J�s��fa@��pj�� ��LF�r��J���������
���.l��4~�~o�oj�.'f��o[��m �r��}Өa���]��i�M�+�m�5i�N�o�,]�ҿ7lJf�xɖm�#���j,/3�$mCW��aLŌ��ٺ�s�«;-Үh���K1��y;_��'Ary~��Z�9w��(L2y� �;�R������#�A�dZ��[���J��8<Z�yEȨ:i�YD�uCM�̑JۿV�������!�?-۠��+�|j������#��by�2�U# nE�8>}l��G -�2;�<�O�����ދ�k�y޸�`:E}� J�o���Q�D�/G3\/:^�n(!s�|dZf��!Ȕ��O�<͞6zp�t��`���tY�ifp8ѫ�w.��O_H�`$�֕�ݗ��Ѵ{��W�f�6�e*���0���	x01��}��L��A���]?���M��]�r��v��7��=�I�O����Kѫ�F>�G��k�u8�ޒ|O���¤y�Vk@��:(���[��߽X̵����[q�`����|�Q�=��B�̣����%�B�!{g<�Ʋ�K�sx�}�T��7+��0�l����&�c������kH���6M���FS����}1p��JU����{c5�/�{`K-Jx�7UΗ�b��Y+Y���)а���Ej����9�χ����~$��������[�����vI�Nqл����-���G�����A#��:�+�"jۥ�H:����>�u�u���>^��J�S4U.T�Tw��H�u�����)��@�s���U5�ľTQKY�»7��	B���a��U�O�sZ"�Q̾�ݕu�����OA��w��%V�:'d������ Eڝ��A]Thh?��j3��VCc�m$l::%1Z�
����z�͛�>��y�ߥS�������u"�.���XY[ψ@o0��:[O���	C��Ȧos���O���[{{sU>.�0����P;j��/b��8�O�lΛЦ`b�~t����T��KH	88��~���]�����۱�����Zv%Ғ[��,��C%s&C�z&'h�WV�	��4�Mi��4�䡢�3����l�=)���8E�7h�#�댩K�M�%\)�Ǎypה��x����2h
~:��m^_�U5J����4�@0B�Z�s;�K���,����YO��R�Oh}�)u
��A��"s�D����z����2[�2�%M��11�;v3��v����!���;Ma,�O+���Ds-�+HW�����ǎc���/�Y~K�P�j8���*��{���\��]ckf٘�R����Kt[6"��m��7?�مA�дr�5D�w�L@Ϻ{�@��HL�ӿs��Df�:$�I-^���E�ʁi'|��fΝ��x�6<�c�4!HmΓ����Et� �0#؉�=Oi{��pc9� �G@�ܗr1,NUT�_ �H��Ҷ�g��<S76���2d ����)S�������^jǮ��	��JFO��Ti\��#u�?����i�X�e���傪4���C>���)�9?y��i����IuN"���5;�I�\gC՜%���Tv{o1��z�}���ޥuQ\��ܜ��^Ä��ܫ¶��[�^
��������F
����ւ�Mo���T��ִ#h�K�w-��Ԝ�]�_5��X�������;�����c��I��8R�I��T;�%x|����Zi�r��:_����GF�K���Tac;�}�f��Ѣ�S���2��c�Ԑ����r�[��Eq8�М�x^�)�e k��l/&[�1ߞ>�q;S��6I�:��B���=�
�8�1�n��OR���x��V�!����X��L���g�HLŕ�wf`�
����ܢY_oҐ9��7�̭��)��S�"���j�W5Z��T��>=V!�3L�j�yg)|H��G(ߧ�g�� ��t[�9j��f��(v�l��#���@����G��P���Z�u�bk��b_pmdZ����mؓ�eT��<�y�mE  �(ݞ�-���I(��z��;Y�ͼl�0��ߺ�䨶f���m�ST�W6���F9���O�Jlџ"����G��,�o�*�w{I%6I�-ˋr�t��� �w���Ξ��>���b�YX0Ͽ�P�	sLy�oT~�]J�MU��	%�p���c�QH��oꋖ� �٫=9�.~G)X*��[p���פc�g0q�ӫ���2���UKz{�U��?���c'� ��]�����@����#���*M��u._�!Y�E �7v��Eg��Sq�F3N7b���"�j2C�?�Ng�x����N��>�coDm��u]�c�̑��ª��ۏ�����u<cj�C�eF��X�U�Bʓ�r��Y2N.���m9��)�`��k�&���M��g�L-@G���n�:��l�L��Kq �'o޴��+Q~:���̺���\�`�	/n ������[���5q���yg�gu>4e�3D�c}���W}�"Qi/y�7Ɂn�����oL��uvUA~���xXv��j�r�O�E�H
󒑺2���Ƴq�����%N�b/�ϰ���+Ըm�ƙIr����d�/�#J��\��y�<Ų�9���O_<��bU�8�G\�|�A���A�2�UW�}o~(�i5��n�]l�d�QIX�ٱ3��� 64_����5��F���:�fpx<��/�U~{ݥ�XO�g]I,|L��r+0����/���u���<�%����4u|�N�_�B5���)m���U��������2��=��#�CӇ�ʢ�����S>S��X��i��rya�8�5�dR�����빋��a��1�r��`���BQ���s�r�@��߈�?a9Nc��=�/�2��G��?�b}��M/iҢ��1���1��IW�~���v�Ɇ!��'�'M��J����$n���q�(tXA�ݡ
�rSx� �c���ټrk�.!d sr#�K�	����aG���QO58�
��..�d�Z3�Q6�7�O���tqyy�";�i���ܴ{��e.42�5J�����	�y�'�T��:���T}���B�Ar��~�}�*��R[�<40���-�H��TD��b)F�o05�
8,�4I��v�6}�^�ym��$%��k�-đ��C��71�ʘ���Td�B�7�S�D�|��B.w����ٿ̗�W���g\B,WeWgbl��������v#
��B��A�������<�2.��+����2us&fD�>;b�3�����('���Dr�=�:'� ��ڟ/��pn��G�i@��gn�<|��� �t�a��n|�k��M�{����e��!���������,���$I�J�o�\�=������0�G���V{��ȏ���{S ���mi�Ju��	>f��Op�o��9#�H5l�,�3:$�wMEkH�^����f,�st1�]6���nު���%񼃲���1�zӷr6Y�oz���| ��g�,�í������)�`���ɔ:EYT�J�_�Fԕ�< ���N\wٱ�R8L��ڙ� <=����O���PQ+RM!�φ���!8��5+���  w�!Xl�	ppq[6�z�;|+��f*�4�_m�1�5�f�8�H��'�z��ܢ�˔��ݷ��E^n�����|ʡ��c̦�,�UJ�.��!�.�;i��$��U/a��&�čl���
�����w��X��0V,��>Y��T�m�"�6m�s�wp�<:�-�R�a�"3hj+Iqi{�����S�0����WV�G*�����вc,��Y��qRU>��X�@Ѡ�j1@�����Tx�,�y��=lb��t��������Eʨ���v�c����.�M����ɾ��q�!	�k�C箃#����!9��c�+�`�{�sc�ʖm��*�[ƙ�L� ����d3}���;���max��p~G�u%cw�o�bi_�Fa�n�3wB���,��o/fM��z����Vz,B��Kv����݌q��]��Jc	�nu�}�nR�6⩘��B�&X�P�_V�{*6�X��rBBЧ����.����!:���jQ���~:[�$�'U须'+���rD�^��?����Մkx�j��G�L\|�L��"*4�|<s��ʒ��ن�g��=���
�»ؼ�W�7�	u+��n3���V�*�Uq��{��YI��|BW�X}sa���}E��,���h|.Hi��YTV�4r���P+�`�`������S��"�SU��qLX�h��NN�0�U<S	x(���{��!�)��6g%e�V���&5�iE�)kŅ��k�C�����/���z�ceS>e�l`Xݞ��oj�d�za��xv.�`��/�I���)%��QҐ���]��:^�ۜ�;"�)3���"Ϛ/�	�݂�Rt����j�az��5|���긽-Qm/���W�#j�C�32*���m�R��^Y/z%f��7��Ѐ�l%s�	p,dR���Bh�~�αu���&���;@�~~l3Pd���w�)[��BDa�E�o�d�/p�#�Q���v�k���v�J���n4E��\��'ʯ��()b�w�k2;����'Ҕ�a�H�ٽ�U�S�r`��4�� �e=l�W[�W%����#�$��U�,��bZ�F\{k�k<vAZ"�y�fT��z/d=� b���*ur2�N�%�:?�/���b�_\:�[p������h9�'��(HU�v� ��L�2P�����؜�a�Oo�CX������U�$b���qj��#�Zo�"�gzJ��?�@�[�~��P]:�<�LN��%e��"�6�Dz�윫�+\F��� ��/^�ڰ��O2������:$p��X�N��O����Po~�V�cc��E�c���`D�J��̿&5�t�!��Ta��E�� =��v��?E.Q��)����l'&!�p�}��(e|�⒪m)���I5w����1
���*�N������Jq$v�.�
0~]��m�;�+�%0�^&�,��3o!�DT9��8��@�"�a�w ��a��1���N'K$Gնb������y�R7\��Tޣ=��b���.{P�����a�T?(^S�~���B��@��K�v��m�u.^�Ǳ������Sc�X���O�宨c�k��V�����K|W��0�u?��ˋK���h�\X�2�2H�!����ꄺxƸ�`�/��a�����&�	Vٝ�.����x����eV[�`.�9J��!��l{���#@��Y%F�N�ʱ��5|���$�>����p s�Q�v���dޓxȣ6��vIL"Փ
��w�ҠWR�<���g��Ţ�| �ŉ��6!����s��TM&����q�ԕ��m�
�ń�L�Z�� AϱT��G �/蚣�hy�]Me
����*�ʱ2���Ǭ�h�i���#??���XU�-V����KV�z�T�r�����~$9ώ=-hf?�[%
i�[l'Ɉ�Ζ:5��'�4�:��u�.���������X����[����E�躬 �D��t�T���xzV�q������}8S��������Ď_�9>����2p5T��10&e���t!�'��xX*j���ʭ�}Ht�2p?�"0L��q�3��ǅ�ͯ7��֡R�;���=t��(�>�=�
>/LC��^���j���(��/���X|9�`x8ˋ7a�g�n��>���	�?/ѭ��Tꮅ�Lz��I7zM�'���m�3�H+X֟���u	����q𑨠+NZEL�F@�b^ޢ����۝iق/f����a��:T�zXw{���\)�s�A;�?��/\zGA��Wj�IJ��DG�|V�T��P����G@�܃�I��4s�z�����h�#@(�5$�a+�}�^��1ۂD�����s��1���=}�?�
"�bOA��xWs33��I��BQ�)�M4m�d
tH�Ч�>~�4A�>i%
سP��հ}|�B
��g��J���y�0+૨R�EH��ȩz^Iw��V��EH*�E	-�[iWf�OLW�<��\���M��YCj�ϞJ���GʔǶ���b�������5Eϱ��x����"��xz���xG��X�#��@�����=��R~Y���pf^ե	�}���F7�hB�N��o��g?�z���|�'V-f�B��ºJ����K�$vk��q�T�fx7��r�u� Q��p�:>�3 ���C��������y��y��2�u��E���\�ХE�JM��IB���O��q��gQ��Z��*/�K�|��T[�[�BTg���g� N9�"���G�c��F���]G����P���q�	p���,��)>�!cl���Ugs%8&����T*�6��`��H�|-��ٚ[Z��Nb�%J��.���L��o3(��-�D������~"2e<��|���Np��!7ڌ������N�k`	�/[�3:w�B�{���/�0V�`�ѻ����ۍm������\���K��������˾!�
��j�H?�-����l!���+N���SS���r����yH�fq7��ܦxs�0�����졭���h2�;@�=���5�O�+�V.RG�ΗfѲ��~ֈcT�_ư�}-ά+��-��-ec.�{���X��'�,,�����o	�~��6��ᣃ.�,���]�aVf �[���Պ4�߇i2>w85�7�/Q��LC���9{��<��.1xy;a	������--3���_�/�Lm��-���^W8|���is���Q�r���qz�Vq�rӕ���_]�Z��k�r�n�9w`���v�<'M��&�~w|/��C舩�Dr�{o��T�M���ewŽ��%Kރ���P��m�s��4�#���V&�%��z����`T�%�K�Fq'k�)�,��S������&���)��5��yӧ�l�Sٚlr4����zZ�b:ț�u�m��yBʰ�bO�peC~�0������
B+���x":la�N�Դ���:l.	��ڔņ����F�j��\�ߞ��=±Mj?�������o�m�M����U�ى���+���QCe�8����ۻ۔Y��&��5�_���JB��:	�웾���#�� 4�|��8N<���m;]�3Q���g������#�ӱu�-���J�8b�Z�a'�-�V��,��S���\���Eh�/4�IUH��-|��}b����#eHL�xܛ�y�w��c�W�e3�"�}O���ܨM���䌣�FD�M*}���13O����z��}���2͏��2�Kc=V����**�x�Au�s ��׌��W�>��k�8X�����)���2~52�?��$�_��q�%�jl�����D�P3�ਸ�a�DH���ް�Vrr�,c	�=t+��{Z�=t��碞�8�N}�?��^Ehw	'�aS�m�U�f��Ig���o<���K^��|�	�<o3)���F�=�pKj�7?^n]'��גfJ~���VlH��Ԩ�$PVÊs�izf%x^]~Go1�v�t��I�W;��E���{	�{�q�ӺTC�3������=/p��V�po���tC��i�F�|��b��1?s���`��g)ٜ�xp�}�	��~X!V�'ʞ��;P���WjU϶��x%��"B�F�)��Lj��'�c�q��1F�?���5�m�׃�_C���t�_��#Oe��[1z���^��~_�$����[G�������k��
�_gF0�Ht��D��O�H�Ox]���&�nK�0�w:`7{�n߈oC��q���n�z'��/���)�{�
e��wߙ:o�+�joSꭚ����6�y���Ə[�o�D��P2�����S�p���=R��^�DiIm�묋�ǿ�:�eb������Q��ph��k�"ܞ���g[���d�bh�!6b����4��8>uV�2j#$v.Dp�t������K���C%�9o�r��c��IAwʫ:�A�Th;�rXi�֩��>���9}x���r���j�'����,ke�ۇ��V?Egvy�R���0����[��r����Ż���������9�e��B��H��]	����jt'�Õ���T�'8�Q
���������~�t�g^�u{�:����~"�b�/�=U��S�@B�g U�y��F/��LCK���5'�:�w���|\˅?$�d5e�����{�'}i�8�Ϥ�����|�@���-��v���9yY �\�o�`�>�P�+~7�˾l)t|G���JY�`Ip?L2��x���c��B^:��W�b�ÈR3�
|�_u7B��RIJ��#���p�z��{�<�_�rp�н�Y�Ϛ�itP��t��F�A��>�2�l�A	���&���r}���QNK0�|fI��>�3��n�L��������>�-j����Lq��dKM5��r����r�D�.�ޫ�����km,xx(���M��k��y�����w��v�|Z����\-�����Ž&�ʌ����D�.�:�������><�p[W�do'4�@:�����b?�5xdD�����y��?��U�7ڙ�)�ھ8%����O]:~���<�~=�=Q���HLڵ�K���P>���S��9B�\I���L�ϛ+��G2��,�2������v\�P�j6����Kۓם�����(�A4�ң��R�����.�M4JGR w�?�.�;K���0TJ��X�T؆p=I~=ޟ�6�1��y�.ʇt��c(��Z`<��M[�&o����=PSY�K�����Qa�O*.�����A^U�.�Ǐ =�/c*�X�(T0�C[%1d�Z��q�>3�G���-K��k�0��ER�8t*�H{c�2+��C\�cަ)�+<���Q	zDU�ց��y^�`��\��V4Q�9$����;�^�ݲ�����Ip��u1���k5��?�XB�
7V
�q�EZ^���,(��)1�@��j ��-�G 9�M|��纛��:
T�7�4�p�����|��$W\4�m��̛�m'�$'� �'���W�=����X�p4�:/!d7m�>�pt����d�Z������:��(B��G���-�o<C�-�u��m⸖���׃c*[����[f7z��M^ϊ@t�L3m�h�yz�o�;�D @fO>��5/Q�.1o�d��lJ#��K�n����瞐fY�g[�r;��Vv�.h��1@����D&(�}̔IϤ۷�f��ɡ���˴o����B+���.��B[F��nmd�!�M�=qU���D�=?�p*���"輯t�\����$yX�r�46����e��W�,���Ah�vϺ!��j	�*\����`�U��b;ؒ�^^���µ���]�'~n}�
d��-���Ȱ����2,xF�ޞ���;�oa����-�8�^'m?S ��0�;�����t�VXΐ�myi�yb�bO�r������co��R��$G-���xC�U��Z!��[�HHfP���z��Z�կ?S38�Y�)[FO����x�GH�������0�58���/CG�ڞ"uF4�[@�~�3.7�, �6�1�	��{���Su�6*���
��o�vJ�qCθio��m�Cu��K���^[I�~�v5�L�������ÞМRE��<���a��xs�p�yy2~) ���A�[�Z+m��!�Ņ#�����\_D�����5R-o�"��ղ��RG�6���rDH���]˾K������թM�D��@AB�z�yF���3ؿb� yD�)�	]M���3���P/�Ƨ;��i{��[/�Dl�9�5��F��Lɸ�jw����@,f����Zr��DXF{r�[%�ъ��F�n�%�����<4��{�H�+�V��W��/���[�"f�~h���0��쌐�+S(/�.�Y	M�a{VbF��T+ wB����ZlN�*Պ���?路ur�P}���8�{o�R�?�l�W��=-�[�ʨ������c�s��	�����G��kM4���m>����
�e'ՌY��mI1VI�nBU��%~�.�|�4��}���r���6�5̀��3+��W)Ӎ]��Bd�)���ʯ�b`N6��*���j�����%�:zbSo+2}���(mM�����`'(�8P���݁��sa�/�~�qQ��g�
�%�(?�;�W���i��Q9��=9 0�e����ׄ\�������eI���ʕ9�l�}�/7�e��?nX�8�Wrأ�m̈́��v�#�d���&��4�~�{R����c�P�ABZ|�����n4ӗK��f�x��:�Ei�\��F��n2Pk[޹>a}OoqdƢ�"��=�Y�t	`dNU�5�K��=�����IA����X�pV9��D^����ʊx�Oй��/[Ftݑ��\˫�^7+���>�"	�=�u��u���;Yl�>�m��jt�W&�f�w��sp��?�8H�![�Y�
*C1E^.����P�3<��!����hڭ�?��..�{���Ư��i�"�i��uҏ��y� ��g���xAi�B�IL%g)c�H�����a�!h�z�M���?3���j��l��K{��������7�o�b`�aa����ʱ4�3r��uH`�\.FK�߿~�x�$�<�Ȱ`��W��2��L���j�QK"7�;�w�.�I�lt�����X�Y,�u��9�ܨM�){������������P����8zC��;�l���t�_j���o�%)?�칻�dxN7�PE�1x�`�m7��~�|7\�_�	�X|k�J�Ս���8ǎM<y��/lL'Ÿ��j�RZ��NTI$���7,���{2��+}�9�b?;^Qv Lw�u���-wA{-ᷰ3y��� =�߿��@*:5��|���[�3�L{�n'�7dFq�:���#I�y��i98%ob�2�W�
d�K�V��=�Wt�bgdU�Mn4#�eIn؆^��jez��?����v5U��s,-U<���J^ށ>�onUz8�e9jX�� gV�f���b]/���f� 0	!ӝ���?vѵt�l���_8�9{�f���E�B
�c� k `�-��hz����{�G �A3�&.��ydj�+�����uI��mx�[�P̢�@\���Z
�B�Q���|q֦��+nm�e�v�
! �#��X�{��h�U z	�h!�	�]�D�w�i����V���3*
��P�XP�J�%w(o$�I�uG��~���n�#�ܔ�`㸔`�Cy&��.�O�z�q[�꧘9�2G��.~�w������+��,bu�n٠�A���H]�X�]��l�_�FcI\�����z��\̢X"z*?I!qA�Cl{����JW��_G:ݫ-w��[��S|�&�>�f��=KG�g��C��I�|���1�J�V6�Z�>�}VHʜ!O@._�o����H�MF���[�b��u�zՍf��Ŷ|f.�o"7Zz?�k�8�+$�<@Z�ĺ~�(��h��HfV^⒠m�qb�J['3YIJo���oҲWX�$�\�f3]�����	f_RB
�C�9���e\����*i=�J�$�c��Q8P����En��f�$��2o"�~%��W���u��u�d�}֐Hrd�ؐ�%�\�X~���ז		�]��bvP��[��k��낶ɯ-���Z����k�^P�P�)�[�_AG��C��7L?�N�Sz�h{Q{�o[�Ѓ��B��a�C{�.�0�J�"�z�$R�J\H`J������E	�@~��2$N������9����ޡ��\DMpa��u�_�,K�$��k^�����F�
���rӹ����P�6A}S��a����S�Ū��*���?��v�Tygw�����Ү�n�I����
������@C���Qb��h����dodNI7l�J]xF��7���11+�`��Z޸eQ��JB�܊c]������
�\M&Xݟ�����?a�aΎ�i�i(��:�=�ؿ�YW ��kH�@���ܰ�2�皬Ց[��K3�����f\���`��1�ɾ���#U�R���.XUcZ�й�����4����׆L��0b��!P��fo�4�g�nd�v���0yRI��g&į!��]1qi�G|���n�����Z{�JwzǢ���ԉR�6j��W���CJ��]����2�q��j���'�� ��[t%_�بP/hx
���Y�<6��؛Wn�u��D�tۜ&9���� ;2;�Y\���o�p"��Q+�ǋ^e��qu�W���O�1m#�r10�'�wG>)[  \�ڻ�mml�e�H�	�|;�UY��¥����-T�K�%�ր+u���y���,�9R�/+��07��.�Q������y?�e�u���a��l��Sy +��9m���|�p�O-&���ά��HX���Ɉ�}�#��1��D��p5�k$�Rl��[@��by�/yʅ/Pm6���]m�S�K�6�苪��7O��vJѦ>x�U�f5�͑��
�SpA;:T���ʿ(�h;4�- �-""0�tww�HJ) �  ��ݩ�PJ�H����O�������9{��:k�w�v��E�M�f�=pg�\jҽ����m�j�
�G�O�{�Ĥ�|�r�,����K�������t]��Z��%�ەy�4:��\Z�:^�-�'�������������v�9���P�F��R�s��^+5R���~�Z��ۛt�˲�mt�h��\.6�tj�J >��U&J-AWn���b����6���E&�RF��!�3m^x��XC��?�&��s2�Dk��*V�5a�b2X-��e�F�� +�Q����yy���x���h���NB5�8��T����D\P^"������	Q����C�t;{�}�G�$��N��M���;^@GFi���%�rO�h�ژehC�4cZ*��o����*}ˬR��#y��}au�Ϩ��ˌ$}�H�CqCXz��O��
eע�k���	�;�myz���?Dy���KmN =��"��`FY��K� �g���(�wNٓn�[텣�H��T�$S�Q+;��#ĜU�ٴ�d:�Clv����Q�KCK��"����t�ܾ�[��W�]����g�2�~���e�b���P�y�C��q������\�՞v�Z�A���׌��$�ku�p!����>�!ܜ�ϧ���8Nb�H�y}?��������g@BB��A��U�������/��G�w��`� �	c^�����yL.������{�T�ByYJ�"\�r��݈%'���u�2ʜ���#̂��~2�S[���iE�!܅R�Y�5��V�F���s|,Iz�"��[���1�iZ�.I.�|Zte��߹�2[����z\�L�=�	u4�|�C
m�|�\�3g
og�����b�6���&�
 !��Bvf�@�^X1�F���m*�Ь��!�w��-ƍQ{7l�)�V_���R�9Mk����Ac~�&�*J,q�i�i�AR�0S@rK����gM���N�'��0���9���c����$V��*{�-�]�*7��T��oN����b�d�|�эj�X�`]��@��4y����K}�M4e�$�
S����~B�Y$�!�E�!E5�Y�}����I���P�*w�в���#��C�{���զ��퉮�]��Xy�*Ǟ�{23a4MG:tT̷1��Rb��kXq�M�a���$���9��zx�Gq6�'����<Ƶ�,���L+9�	.[��u�ʝ_u�x_����`m�iK%��ի! ߴ�Pr�43 >4��噰� �(N�sX��S���r��E.x�'S���E����o����IY�(��i��sɳ�:'��2j�㒕X+�.�R����%����V*��x�"�NJ<��Ņx\9rN��HT�5���v_C��N�;f��f�ĕh�����ߒY���$ȟ@&&"E?��<X9j��$�h��^�/ao&G-l��]nH����7|&Y?�D=�f�^��q��OJ����ǴV�?"�@�Q~ͣ?-�>��I�힄���ER@�T-C�o������&	�/�k���o��ՄVrYV^���9�~�s��ת�HG��7�X;ۚ��y�/B��W�U
 ����f�����$Hᱤr�A<��P�}�S��c׶��N�����T�a��\w�˦	'�*>k�Ę����V!YH'��c���_�B�dx��?�뙏3�*׌l}+���.�61L郔X::""~�:)�7�3���(�@�õ����Ս�ʱx���?��!s�K{bd"gf
�H��δQ��nY��kl@?n��)���m���0�G~�X�WÅ�9���R�>{�����+�F��?��V67�&ק}�Q���i+�eF韂f_~ؔB]8���!����?3���������=2��:)N۫O~�1� ��5��Sa�nE��Z�hp[lfT��͔�tN�z�2��s�f�t<�E�k�"5"..������C�3n~�Ҩ�ƫg =�̀?�Z�r�����F�x�*7�(/����e�~����tp�4��W��^�?<�o�biq-ƒ�X��˨v�W��Ml�x���JVx�uSY�����x-�=����S�q� �{3_�1�P��AC��^N���$3\��@0<V9��6��A��hPO͍���H0�`��%
�e�[FUY7͐js
���x�2`�3����B��^��b�lXV�� �i��4��\�	$:Jh��{ox��F��;W�ȥ$_
>����R�,����6�7��)����W��o����#�&�c�o��H��\\�چ7R��m��>N �O� �g���ߵiTf=G��f ��O������ѐO�Vp;���:ִz@|�T��������S֧�]�����g �u��]���0���J������;���#��VN1ڑ�w���佚P]��7�$��Ү�E�-�� ��߽��G�������Fhq��/#����0�_��K7ֿN�[�(y�����2>�V�dd��h	��۽j
UX��'��*1Ǐ!���.�5T����~w�- %_����e@�u/��������x��kd0�8{|,�^Q���E��[䎂:Ԭ���e1Z�<�^��D��Ѹ�_"M��E�I׽���I.���R"��1��<_�
�W�	Rx�x����qG�rbHm#��`�~��*Y�U@���ұ�00�D�豥ͪK�R�}��]�AF�3�{�5%��O�0"N�{xR��{�#3$�<�h7ׄ�� �r����Э����`�� �o#%6��2�;2���O )l紩CK�r72� ����j�=��<���(4�k���7pd�I*��9����6U+��	%*;J�ȿ+��}xs�x���Q3�M��&����b**צ�pQ2�m�tG���$��,�"�;�6I�H�������Z9�D�g��N�>������:�5�%1��%&SI��ysu=�#k��~M����zn�ӮU0�9���0�.UF���ϼ���(9Us AV�I�N�ʙ�Q3,˩OXt;�š��y��1�M�ނU&���Yk'�s�=x-��W�2��lI�n���bj�F־6��O'=w�LJ)����No߯�����R�����*�1���;фi���ɺi�$�U�;;�D���RM7����ZD� 	��&!�H�h����DMq�
�[5'���x��uH	s���Z��J��7�<���1��c��&V?�7M��է= �\��}�A�� �wY��^�1D�����
��X��%$��<��K�p���F��&UU�X�Hd�Ǯ�����I��˕����N�[_h���Sat�e!ԣ�MP�T���
�|�_��W;>SSϣ=��j(�w}U��3��g�Jݿ�1��x��S��eIҞ�z��Y�NaC�V_�h�M�t5� HS�D��F�]j}}� �������l��l���n�k�xkJ��+\���{��I}�^]�8ϗ�5S��թ��b�6�����1��<���q��������.�!�j�8)�|,̇w����6,H���'f��πJ$w��J�=O
j�5p��I��@��!
�#�ـ#c(��m�u3�c�S����/"����ZqRLqg�(]f@G�X��}X~˕�U���Zk~I�Ϸ�k0�═A��G��q����z��HPS+�W%���Z�č���}'h)��VD� Z!�5��Eg�AN�$�h&s	B��f)r A�90��Vs#݊�W��"��9$��,	=<�bb�P������j������3�z��8b��,�5��F��,�kJ��H�_���*ƿ4�gNp �M�u��J�r��kBѩ��_�z�6d��&�_sI��bT�f���Qd,������v�PR�rc¼b�����tq�L`-h��(%!���o�۞��n��>�Z�4s�A�����{%K���Q  G���3�ݰ��k�d-����r����
�������P �|���-2S���nG�y��|#13�Q��7�,g�?N=��ÿ��+Z���_rҘf܊:-�MaY.��z�n���B��g~π����:�'�#�1���&�v��Ko�y��-��w��Hڮ�Iu󦆸��=��%2n��F?���4H6u�m(��k?�"������ת�]���%��)e�Up`�p��8:H�����R�X�>۩Ct�ؿH.�bORK�Z�d�f�wܕc{Ȝ��D��9��
09�O"A�L�dS��|��!R��_t����M�π�@
�u��Һ��2�M�uC#��nilQ���ie
O��i���OX�KU1=��r�q9<���Y4�ی�l5;{���.E~	_���q�G�8�~���x��P�,mBzN����]�hHy]��x�2��^��7��
�唹0E8Q���7a��:���[�s^���k���P6��].Q����ju��ʮ84�ֽ"F�F"� k�JH;D���*�ի�֫�r�RW���0���g2�R��?u|������s2�P9�}�T2�X\)Y��)�Y!td�y�F�Q���6K{�iy��o�>�����j ��F���#p�ywn�~6���c�Ҽ:q��A~�^]]T^�*�1Pjo�zI����묮��{#��4e`�����χ�5���1���yFƹdꅶ��ܺ�����&B�r�{�9E� >zk�\"���2}���/]����Unx�lKC�N-����Õ6��N>Ť�,�#�(��	'g�u���j���6���au�a_��uS=:��rT��@(qb3�B8��*S��W�9{t5ۉ�q��Ԝ�P��٦u����1�}�NNK4�bu]M���$._����m�B%��>QP"Y�5�c���d��vZ�=�J���-�3�-�H��_�^?����1.UO-��k�y�1��+HZ�?�K{�Ih?�(���3�%�t�=���OǨ���%�Mv�׈ �x9�Q�ai�mC�Rx�~�%��Q��/q�>���ìW��8��씾�m��H����󴫻��f��/#I�	I��rl|2?7��ɘ���hz˕Cj��:\�	<�?M{G'ޗ�E.3r�����?��2��˝r�$�9��~,o�R��b�;�jڕƐ�W�x�'�WR�IY������O�re�^��O֡��>��%9~�c?�8 �������-;Ys�Gq���R)�ia3�"�N�c�䶨��p�AE7��<\c��J�����ƿx�/j�%N��U�,�9ˑ��ދ�Y�G
4_���a�PX�˳�ߪ��)3P�޸��^����L=��R�r
��\����L�mYs���捚�(QM_TA�__Z^���w��0X�` D����w��H�1����	Ws�m�5A.�����Z��8c�U�Ή�J))�G��J�uCaL;V�'s�g@���8�w$�J�i"/Wx��B��8���9¾��֧"��j�c�P�iJq7-C���c}OTK���c��f2}��BY[M��*�f�D1��a �d�!%�����DCo��'�v��d��(ԏ�u%
��|��	�7��0�C���ͣ��!u���/��˖_k�M:S�����J,	�¡&��6�3Iƨ�텎Cr�|���)p-��%M}6��	��d?!A�D��k�4��:���6�� ��/�S4�}�.���t ���>����w��ǖԺ�¥/�?Cux������ۋ��
���GA�݆��B$�(��sw��4g٭U���j��K7�����U2L�ଋ���5�ǯ���Z��5D��1��i����U����C]p6_W8�0�G)����b�?� �F��r�>�~sr˩0AR
e{��gO��E�u�x�Zh\���'�	��(rpP�6�f����2)w��_���]�ښa~��q]�A�Z�o����0v'����z��|��]��}�m:}��I�����<'�۳VWB>�8-�;\�S�x�4dK��J���e��3�����ة6��/�.�D1f����'�O�]pg��/tMA{Js�]���|�z��9Λ,[6��a��dpq�ٰg��f	W�};�r�F�`@�L�}��kӜ�h2������h��T�!S��f5��˺������M���Y�g�d'�]X���X��6��ժ63FQd��<���Pgy���V��~C wy��{+���g�?�u�dt�h���i���IW���Wt��/J("�@���,��!���a��&�N�����Y�ʮ+j�?��M�Hݘ��/!��?���n_�L*Vn���j�gp��7��o7ү��B���m���!��z�x8�%J]]����d�F��n��#��uPv8�ʾ|�������*K��l���밝�-x�-�qG2�+"�ix�a���&���'8Ew����Zĥ�U�Ո �]�˚_�o���䦴���#T��L��r��"�^/qp�AC4�[l�~�L�7v�ʏ)F�JK��.�Mol�6"�k�uq�cC�\�B:�B�bV���+l)��~3c���\���=��Jm��U�WL+�j��'z�$��SĢ�>��ג��CCfEF⑥+;)���?����l��G�I�ċ��LY�Z_��x���巬�U[1{�9�KG���M2��H��4J�T>���*��.ygr[�o��ߜ�e�VH���Hy�j��d�iL�����w�M�\�~��=P��/�ȭ�K�w�@և���c���l�����0SL��������a\8ɮ�w*[w1�z4�6�]��|7G?��{;k���mxb���8aR��Z�W�z�������-sc}��	[5y�ܪ_�:��(�g}�ۚ��^+e^ ��s܎�0\�����Mw
2��i�G��#���F"���u5�G>�]H�ǯ'�9��e����V;+�
v�+�rwr�)��A�8�!���[O��ʊ��)�]�7έK���>]<�W�Z�wB%��.wA4{T���<h8�J
�PYp|�� ����;_�b]����=���XcЄ�/Ô_�?0��JY��'w�0���J�y�?6&E$	�����40��h��a�;�����i�%0�k�:kd����2Ŕ�����)��`��']0��P���t:�*;������F��ԻEh�XJ��/_��""�u`cÐ����&&���Xx��Ĭ��%��� ��l���Pj2<�����.��2k��lJ=��cc�ݓ��C�\i��3�������<�R��7ת�dMW�.����7���_}(.j���v+�*
K5L(b�V�~	ȽZ.y������ณ|���x�x����%7N�ʪFMA���B�S�P���~��8��oy@{�V�6{>���׻�C�	v�j�����d��4c��4[oj�?Β(���?v��~1ґ@���q�b���*�ϗo�٦��oz�X��Z��rZ�\��v<�e�w�[L,��T4�'��ݨNAih�S�4Lc���2���g���b��E�O�0��x���p�z��[w�a·���#[��w��i ��� 2�MU��p����,�k��Wi��N� �8��~��_?qG����V�.�V�o;�9I�x�v�ՓY�Y0].e3S�\����nN9)�%�^���o�����@�g(+���w5������Z�[�_��#{Kh�:>_[<����w��W�WI���B����S�hsl���u�%.�d9H��R�z�C���^O�.:�M���H:����y��v�{��������I/pRpI��j,�0����]��� �g�n:l�Z�. �� H�-;N\��C��K��ՀL	2�o#.w������ܠ�wB�D�ҙ>�r����=壡�d�h�WX#c��הha!X�-�� �/�~�� 
9_�ƝS1Y�v���8���"��A��??zew8%t��~gn����\(��]Xs�B�I��⑀!�W-��X�4T�$�6%h�����;ANj�g��UI��Y��5:����C֖�zu�4����b�h���z!�%���%�#�i��c������"�7��_x%e���@75��*�J����5I d��xz:�3�����
��o��%@��n����ԧ�}�ow�������E���N��R꠱�O�D\ ���L���}������ؗF>V$�1�������衪�=�EGfz��|�T��>l}j;�����24���eĞ'�H?����I<��G��g�_�. �9�fP|�t-D�<���� X`��~�(�3�Z�az&��j|��h	�O�#�
f2^�R�V*b�(`�Gh��� ��-w=c���&Ҭa��J�����T���2Ny���c���Q�U��Z�؅Fr��%���Cz�ʰ[�U�9�+�9�w7s�Ki����G�&���ŋ����||���j��$��� �ߔ�Z=A�n��Ƥ� �]�X+Y��i �y�
Z�֋��_[�*q �|�A�ng���xDM숆���b�f5-O+�bR$|��vvӯ̣	!}2�/I.����O�|=?�h�U%�JAK*&Y��~��o�٨�^
2�oO�=}�v����0��4Մ�l.�Z�Ʃ�<�,�??�Ϣ 	�QM���s+���� �!חWp�,m(\�1�;���3��ޗ7��S��lgY�EZ�������LM1Ũq���G}��Ay3�����/j����M���!�2��
�pY�۹�f�`��Ap���)���?Kw��^P��.q��:��˴W
����b�:�֫��.j
Dpx��V�a�D���?�4���������� �����v ,k��.&s�7���6��Ci��qj�d)����������u���2�x�]>����A5�ʷ�~8�d;Q�ߥ�8��&:ھ�ȷ��_�f��~��k�5em2���ʐh��z�eINU}�,�!k��I�����e�[
����U����$~���O/n"����*w�����ܜ̬�-oB��O�p�C�.�{#���c+:��i�o�L_�dϐO(���Έ77�(��b�e�C��3i���D��p0���ʔly������P-Zb�VH��"��ځ����x�E?zHd��>� K��7H(؄�V�0w���&�k�Tt�@'����~K���~~9d�c�s�xMGn �N^����(� 7z�3����ލԽK���Sc˴���Z34�{I���S�����4���9}u�$�OߖHnó�|x����K-W�9ü1�Pd�)
d��~򮫥�+��=_R��*�9�7�
��)�+��#���/��S��)���w���;�(����x��-��\��"�%:�JY_�-������(����Ίڦ���b9`������W~>���$��ƙ��_����MN��i�=�ң쫉�1�?a#d^�6\?��{||n�λES�n��f��Z~M�|�C���(�y�۠�������P���L/�^�8j~��$���*SS�4�Z�:�ڌ:��|��iھ�4�H�5��(.^��M>�6���)�JQ�e
����*�iYr�j�@��m�d�I)~,p���V`v|5ǣ�Z�^n<)+@�|�$��@�����zoc u�~�L�(-,�M>���3���<�S���z�K����mWY�oZ�pz��a�&M��´Mҷ�H��x��H�{���^�����������'��)K�
�F������]��/�����mA$7|�TƅnN����0�2�̲˭���[�W>M���;)�K�Ǯ�=:Ob�����l�gy#�~�ů�����^�LZ綪�&{�T����Ԧ��$�p�k�m�J�^��@HM�FM�f����Z�]�Z�.&G#N�~��j/g�k�kY��,��H�|��j�q^a_:-�je�&d�������A���R<�g8�_n��D©C�m�#�>'*���>�.������]�jB��U�v��T�j|5@��i�􋫦�\2��������/�5�sr��r�}%�s��`�g ��X�Iߛ���ݨ�8	e/\��.����1�&�ݭn���	��(�GYx+����L�3��k8|��ݟ�U�:�IЄ�(^0����2�P
����q�|�X��Zz#�v.�����g@fQ�v�C0e�ߎ0�k; |����v7�L`t?
\���-�����
�#AF�^{�s��D#��_�X:�Q�Q�Z<�6Wq�k�>|����'�eIIș��6p�@�R�����������j����O�{�+���F��C�F��B����HS�z�<3�+�FT5��,���IR6�,HT�Q�dhŒO)+C
����0���������ǭ� 0m��⢊�j�a���-}�U^iN.�I5�����tK�E۸,I�ڙ*޵�?�L8vp�j��!)�, ��`^���A�֌�$���n(h?�4�g+a��/W岪���%ʴ�ȿ���P�W}M��@�w��Y��ڗ�cU� �>�_�=����ԕ�Ni���m2�#�IyJ��bXӪ��1tFt���%�c]Ә�@��+�-���?i`�Zf���4W�J�z�i�6�/z=�=vX<x��~MQ蒄3��a�r��WS�a
�ړ��K���:� ��O��	>s1�9�&��W+�3_L"�fi�x���!�_1 �r&Ǭ��6�5�{�hS�i�t�����fvB҃��LJ�\:���Z�~ �B(��%����)�e{�Ҳ�2���B��MM�L�D��d�0/�|ұ����m��:��s\(bJ����*��e@��懕�s����[-U��/J�<�?��<��?-A|_��i�Úި�e�7�ޢ���MAU�8)�IU0�
J��j���ӌ��^�$/��E��/��7�cy�ȖSn�.��9pi��#�`���o�/�"?*����Ѻ��&��p��,�rN��߇�.����	�1��o#��B0/p��g�ϦC�ɱ�S�h��G>�׺ﰼİ�w�q��&h���Qx����7I0�)����}�}<|�OMk�,�6��Y�4ľ�Xk���_lNΫ���%��L�Q��k`ʅ}4���R�/^hnVR���؆BF�$����y����In_Q��ŕ@BR?�ʗ���O4�݉{�&I5���sž�։Y����)�x#�֜���ՠDP:e	�s*��S�ȴ��^yq�`KȖҷh!���`_o��Zajs��� =�V�*Z7��ES��r�֎����״z*���#��*����4.UF�Bmy��o��)L��k���o��&�NV���9������T^�� 
.�}�a�E2逗w �o�j��ffur��#�[�[�F�Z�8��R��b��߄A�OT��+�p0'=���*?U �C�>�6��������Bw��}�(���Q�kUb��/��(K6����C���ȧ��i[�T"�$^� q�X��|_<��o��M✤[�0�:���f��;�39ñs݆JI*�D������i*Y�?UNi�L���u��,o�g�O���I�sC����N�R�C�6�F1�R����H/���s🽃�#�O�Ԓ�X�S�I��:�W �'��[|4�n�����`��c5`�y�� tF�Fq/�/P����k���W���F2�SelL+6%��[��џ�p�X��iǽ:�NG7��ܑd�((��K�J*�����`���6�6�@�A�};P�-��,ܲ��>}�0y].Ş8|&>�����#h��w�\/`?4����>��u��8Ŵ{%�.ݨ��bH���j��7��{��{�Ė9?$��R<m�Sс_<��k����$�E���@�C�% l��!�� =9�^4��\���tG�%$�?߭��?riw�Ya�|7�SLD\:��db� Z.3��V),�Aٛ�C�:�֕8E��,����D��s>��|3�qMך�Dg�.2�힠��/���c׎g���@��@}x�O�f��%K��� 7���.��4��%�pW��v��'�?R�����������t����JL^Ӌ��Iw��D���{/�v��jm�}���9r��iW�	r�0���n�w�������2:][����
��=u�[��H�ݙ�/
�Vp�i��W|g4�����'#XA�/|�%ʹ"eg����]�@�D�{�;�*x���Hxt�`�;`��O;y2�g>�W��x��+Q{t��)���p�w3ÿ�/O��zE`�O�,�EF���"��N���mkI5���Q���A��yG���Ֆݗ�^��E�K�L�/t)�TUA��6X1`�����q���;�����xw��A�-��|�B떕�0Nj'@hF5�q��C݉���qK�O��-9#��B�4����x������o��~>�3�L�Gmd�܍��3���Ngo�-���[^6mXZ�{GY�7�����m�2;��Y�H�#��rHf�ŽZ3o����l��6:�K~Y�W�1��a\lp�!�</����	ua�I�난�8n�W��>�{���%z�dH�4�(��`ˡ��a�'T��bA��O�v�Q��H�y���',���3@xf��Q������4��~�}�#��zP
�Lc�P�n��j�آJSk���
7�b��b�^����]��&1>V	p\t��ae�g���j\q�`<~�)�|Y��[�'��u)����`���m��Z=W\T�z{VC���Q�Iѻj��ȘoZHM�������� �=(ֳn�-p��%_���פq9�����u��05xRH�j2؝�p�2��?��я��ǽ���:7�>0.�snp�e�T�N��t�P�CR�I�ןi
�_�C�qi� ��B��\'�/AK{h~�tS�;ː?���Ȑ9���YkCQ�3o���6SW5C/�kC�u5�	y򬫋�A'	�G5?OTO��D�l\�W�/u�j�}.b�j�,*�]�&7�K��e\S��w5�rbcp����Vuu�L'
��a�c%ܗ0�6pJB�1c,$�5Z��G�6]��-7;>Z����5���u�g��ʑ��+l��w|:��d�Z|CQ�f�g�z�	Y�̌Ua�j績��f� ���I)�Z:�%���M����!�	���G_LEaQ�6�#�^Xc��I@�,�$�`O�?>v|����x���Ȯ
KqR��<�b&	�~kl,�D�xY����Ұla �Z��V���kE[T�^a��"qܗZ��Iэ���?s���VU�?�nl��;�̍/桬�������.2T�mE��e��̓5{}R�{�k�
���� ъr	Uj���t������I�~N�}��kF1b�	㿇���[�y���*/��=|'���b�TQ�|��f�S�nY��Y�^���맵����:f���n�Yֱ�n��h#߬�v^���I<����,V�p+�%�������Z��[�T.�7�S�,��[�ny�?UO|k�~qB��,��z��:���;ye��/�i�yܹ��X�}V;��;�أ���g�'���?�N/�ק\l����X�r\�fmV}zq�w�.��#a�'8�6'���-�|U���,t��������N5�n�Q���%�Q�[ �ǩ���|������/�l�_��_	+S�G�C�P
~�x�=xF8֑��0k`
�3'��8`Z������ 6ߩ�����	��"����J��U�H��i�����n��ʏ.|��R�����(!�cP��4�+��C�4���5�I������a���zw�#��?]��E�Y�Hl|҅�$�~4��6W2�h��ii�z
���n�T%�@$���� I��9���ȏ��I�^�藶l7[���6��D�4�ʂP�W��_u�o_]�P(��A ���P�SY|�> ������qC����[�8v�Y����ɩu�{��~ҦW���<���TA6ݻ#FX�<�8�ȂM��S,�� a�|��Z�9)�%��I	vx5����O��^k�0x��^

�2ƒ ��#�4��o�f�� X�o�o@�[{V��M�䪥u�Y�ǵu��o�xr@�N��E:9;Y�o0�)��R��8c���B5og�� ֟??9�>)(0����
r�*��A�7��_>��ec|Y�j�|���������<=��PZ�\0u���XJۢ�9'B�Fh],L�$���ʫ[�p�H�i~����	�b�I��	öfuU���/�7��7�g�H�4;#��`�$��Y��bp
�zѪ.c8����� fE���׀��	���5BC���:G�Ὶ#`r�z-�b�g�_����D�?D�:�^<�u+Bl ��P��$�L�{�i�Ot�C����w��WBb����p�kNa
�|Z���kT����WV�(�5��f٪� �ZB5 �����CiQ��X/���!L�p]\۩��4�o��{7�yDpE^�B�tA'�U�w�:7����`����)���Y�1����y*nN>�z�����彡^���Ay��}[AVEǵz����d�����0��Rk#!.����'�z��8����î�����I�VJ����,��7_��<�B��g 䪜����+��3��jcSL��С'T��eBm��~��a���r���ʉ��h�O�חޘ���-����cA�{@8t9�S����]d��t9�t��w��U�O���n�*��c�����!Y�b4Z���-`�~`�d>�0M+�^	����!��(72�2![`��P*.����Ԣ�3�=��;�pm���fR�����ğ�r)�%ay�Wr�0l:�e�_��Z��HXL�(T��.l��p^�t�������}_�'4^4T�7����oM�+�)(��JڜL��3�q����-�n���>�ݶbн:��x!��w8 ����� ;�P�G���KI,F�$���K��5on�8����x9z��oW����g���M��AX ��B��Б!�N#��O՚/�M�����?��X#x���َ�:�ǁE��~uee�LtFU���I�]sD��e����l�{% U�Qq'�A؛?�,�[?M���ìZ<qa�=4��gѪ/y)�zo[~)$��"Ԕ*�������*F͜B���7&�Q����=�O�e��)1A�,P���\3�.�ӥ,e�w�M���Rg#|��;��|�7�{�UdNwZ���`PY�����5og�48yҮ�@*�*L��Zޜ�΋=!�Ay�6�B����߱/7��k����Z�\��3�G}���:��qHf����/9"%�UcF{J����o���?~Y���U�>[Nh}�>��bcij�%��m� _[�<�/g��MWr%?�ޏ ���Ֆ�eÀ�d6�t��e���"r�r��xaW�cH�F�Fp~o�$��<:̪o�;%7}��m�録�a[t=í�*�'�Ҕ2I�j�5)�;코x����{�����Ж=�3�*���".|^������5o	��G��aL��%����R�#sg�o����Q�o2P�E`��pO�/,��l���BV4M�75�I�s¡�����|��ƃ�|�**���Arq�eB��}�o;�gc�U�y�� j-IG�=�M��GZ�Y�/a���t�����4�m���9j�\������R�X+H~�)�X�/� ��okA�w^z}0�S)uc������厈��&���zkEL� �W�Fǒ@I���"qGi�upe����C�q	���o�4ũR��2�)�5�(��+2����%��)y-,�,�h�Gǩu�m�l3%���q�x��%�ҥ?��!��~54�uNœ4zQ�E�P���q`X7�!��k��f�akw9V���\Jqja�ib�h��2�ҝ�����kg��nZ�>�م���eo��#cu�L��Ӆ@G�uݑ��/Jr���Z�T_����g��;������p�����r�[�EdU���!;b�n(%�+e���ŋ��4O�nÛO�7��%?=�`�$��2��!��8��S�40�Q���_%L�=m��������쌼���y�F�׿'
A>����leX	w�,�6�\"�������a>񃴊F�?J��9ޑ���X0_�g �h���}��x�����"���
��B�g�پa�/���A��
fC�*��������`_�ȷ��jY�0UZq��<�T(�Ef�K�~�vb��AQ*�iIL��I�AU	�ʚ��s�z6���?̝�CTo�ǗF��C�ZB`ɥA�K�C@�[Xz�n$�K@ZR�AX���O����WϜg���93"�v�_p}u�~=_VQ�SR����RQm:Et]gA*¡�i�Z=-���Sb����C��-�"���F5��__��V��Y:�;�����D?�T*bj�;!/���t�������jfM�/���}j�$>/ػ����:�8��4x/|�R�TXf��f�vl�]zl��'*9�[�ˑ�k�N'�X�H:��jq��7ю�tsC��1{QsG�t�Ȱ��	�²��I��lڇtF:��rd��>"H9Bww�zo���(���[苎�������4D� �xO�l��+�r�Q�!$��"���
�	��7B[�v���0q��fs}�9}7�q��F�3#�S���N�Q��x��
��3W0���K�� ZWM��_U��	�J��s��K�#ʰ�������B��Hz/�����L����)\�
��/��>1+(fr<����8�W�����e_�7I��\RN\�c�Qǰ��Mܟx�X~E�Pi�l-��n̋�P�����#�7�B���C�~�����p�92�2�caux��lJ��g�������`����sϠ�����r�v�Q{Q{���'U�|GFjXi[���/�-�w%Y�p��S�����]^��	r�m0w�¥�\�g�@���C?��J�_�qk+����=L�Z�cL��8��+�9�=�h n9x6kBN-��f{�#ڢ��Ŀ_i�)k�~t*AR����c��8Y��}�[��5�F~�k�DK.��C��1�Ǵ,� H�!
d�hEBr?�7`��{y(�yC$;!�����QGE/�~M���������$�]�E��!� Zok$`*��9����YK54�C��^P���9�&�V�;�8�*h\3�m�����I��`U����1`Q�q�`��V��,������2���K��G��	Ne�g6��0yqrp@� �4v(1����J�2�w j��M�����I؟��Or�v�;�Kǫ��LF�.p}�ML��~�v�
X�!.Q ѯ�/\:c�i,`�I��nw��7�s��nH��'���)�p c=8��C9�q��uFꈸB��_VgPW�ޓaK�NGQ�g^_���R���<'�qR5�s���e��C���(�����^}�>��;1-�bڳ�Ol��LD�W�{z��{н3�W�Yџ�`��mQT����� ��w�j��W@�!��	{^�j
i���Z�eqˆE��	(I�t�:�TW? �J� 3u�J�|W�?�'�;;6�7!��S��A� ��al�Q������e'p�N|-,ˍ()CG�r��10��!�~�Jlq9�o�3�� ���t1�η�M���͕�{.~�e�Y�7��&�o�q���85�E�������d�����}���ҋ8�ip0?n��$��m*ѡ��������:d�zLAN/����d�����ҕ:��hL��vq��O�[sÊ��9?�#_�T;,໹���o2�9/���9�#;3}%d��V�O�RO��h�{�:=��؎�f��A��i��b_p��������'N�{?cQ�Fm>��K�`9�Ѷ��	֘���y1��L��'Q�WI�!���_)`�}��pE�� �w-0P&�� ^
�5�i;�Xԇٮ��?�C�#��D Y��̹�r�`<�D���-�$�й�\9�!�@6x��!ڕ��	�X���=nʪ�jxݺG����%���۔b��䅾#&M�;�@�Y:i�Os�d|��JS�|�?1����9Sߥ���z�6/$`��n�%�j�)��� ��h]:��w���z�] �u,�ƚ�R9 �~�Q��
c�G��}Az�i҉��YyL]�Vx��x~��%XG1�]��Bl3��\l�����ți�z�k'#;���S�qj>͡:�>�f���,W�'���?r��/|F��i��xQ�z|զ��4#�N�YZ:�����M��vxX���ʆ�=Uf����hk�1ԐѠ�|����e�pӦ��$D�rr�xK+�jOe�W�\r���O�\b����RF�Q�t~(��3%}\���ac�h;n���ml4g�o�M4}�4kH_�������w�=�t���<��K2�D��D����==�G�Cg�(&N*��A7T��oG�C�g�޳��Ҧ��)h��>nׇ���C@��(-�%�Q�T������Y�M�7=��<o�����n�b �"Y�8����p��DG����Mc+E�[�?���{����2o�y0��$�;}�������J���DX�xX�x�aii������A d�-�=`B�Bk�'��0�A�e2�Zp��bo��1Ǵ�ryj��PONO�KM����M�؊�������3��MK�{��D�$���S���3@�����c���7p�S3Z��C�L��m�ow��>��Q��	;����)3i�����e������O�@��j9u���'	���?�����{�mK�����fvS��h<_��>��`��Տ��4iG�fzJ#��MZ��Y��=��Gp���2�z�x��9=�W1��=�o�A X�h�}����X繲�&#��1"�+ ��P.JK i1�\�-��MbXm��H�^�sT��tw�,�D}�	�uV
� Ƒ�a�쮺���j<�u�J���iP�c3(4�m�wvq��N��U�ݟ+o�p�D[�h@@^Lz��XTy"��w9�9r�.՘�A=�fU�C�v�Z@յX��[��������L]`j3�Q�� ���D��,g��2�<��Y&4^J#\�H]x_�=�yT֘�s�`�$�d���;�JF�9�,-5�p����?'��d�Gp��ը~�>���r7����B�~C[}��$!��.��6o�����\��ڔD<�DƅEr�U���\�F1��L�l���V)g��Ԁ��G��څ�s7�`p�s�����c�0B��At�2ʢn�l3��^�a��cess����W#��l���8�=b���AU�/�K �hF 4-����1c�Tͩn2������~�>(�� �Ou�	&Q��v�&�'%.�����# ����e�Y�b��itv�t~{�&	�$��@�%"����I��8?�������0,Ǽ�=x��k�&�ax&1�U�*Zk�bj@Pm��=��Nl��>�W����� 	\K�N_��8�7G���b�%�8�tw�(k��q�㐽�!��^c��\bY3՟7)�`d^� �_S�)�䡱P�N�)`���Cm�n��h@�bbJr9F��\�s/�q�$j��g9��މ�c�J�R��2Q.���%C[�Ƙ�yh�j��r�٥�����j�,G�c�Ki]i8f���9���K��y�\9M���!�4%}�9P�� ���9a?݆���7�"\I���V�oyǳ7�ӂom���:����A��~��o�-3�b�b �������WƍY���?*ں�xq��w�;^5FP/X	�x��U]�V���b6������r��-���^b�"c%"8Q��y���WӋ�9���=>��+���. �
��c�z�.���(��M�_��:H>�]����{�+2' �2}{4�u1~5�Ӈɰ/Z�O�B#�S���c���_�_Ŀl�--����\v�\��O�k���/D��.cV������)M���h'�o��u|"Q�K�/�c���e�������)�U�۠�
B���(�-N�fA{2^�E���) �Hm��9���銄h��y��m���g���@N�!�574&��ۖ�gA��.�Fخ^���ġv�*��G
uq�32j�1|�|��è���>�&*�bB~&^�KL�5&��DˏI��ІS�d��L��#�IU8�4���n03��?ȥ�����k!!�dPm��(I��� 3U����ln�H�f3� �:)����1ʇt��+�G#�|��w��뛓xc~]m��*Q:���=�H2�O$-e�5��7Lˈ���i'��>y����ۗ���+cN����SbbyE`c��<N>�W��V�;߃N�λ��I�"��[�ˁ3�e��9;?,tѷx
���>����|��t0�B�W����΢�<�%�r:c������aY+��us��Y~.��_
�U��C�l��L	�&:E�J�
팰X�ҿ?���,�i��1qZ�~��6��s��LH����N��4b���9�
��y��'W�U�p�\�X���%�zL�OP��-�NU��� 3�Xr[NVW�K�e��_�q�\'��`�6Ft��~�����KHhwEN�S���ܾ�������=
ǒ�j\�AN���O���c۹�^>���ɧ�qC���"�5�[���%?��	S����̺;�6^�EѮ�s��N��zZ:�IC֬���+�ߝ� �����v'������v�TD�;k�͚L�j��i&�<S��g�*�Z �����t\�����B�{���Q�:{88���50/	s������z�ퟚUzC�z�(��Bnr̧��T���y�:] 0�.Gym������3��gg�U3gkotH�-�.�a�YVVho���ɻ]���<TXx�Q	�v������n�?@f��V�����!��s%�tXX~1�nЙ�?�h�c���,y&v?�0N�(I�����'~K��F\�1��O�C�N����e˃�n��c��܉��v:��+ W�C�*k*r�/�]ax��`��������R��� i�G�m���۝}d���!(�=ZlZ�~��D�m���v{璱	Ep�]w�M3�@�<��{�uG����ze���g�oXk���s��q��\�ص����ufW|� ��J��'e:���j�D���N��y��I��J2��z�&Oa�ޒDFU9����X�,�7d
�h����ʊ��a�q^�O��-\U%�G�y�{���.(�7f��d
�|�poj�ɷE�\���W�Ai�.U��#����E]a^����� ��?`K�Uq(Xu0nX]�����DY�(���./g�W�͒�<dlq�9�c�c#�ғ��ec�Qq�?�u��!����=�����w�yً_����f$l�J,^L'*�8*��ѼD=S(�>���#m�X��u*�Ҟ(�{p�[y�ڢ1J߆�\�^(�P/�����#�ez�W
±E0xLGM��&��u�v�C�q�r��\��sś�0�.L/��E�"���[#V,�3T%���'�ys�4���s»p ��X�3G�	�0)�`{t���i;( 1~(�AW�+$�Z7p�>]���R�MY�\�7m����Q����q�nl��e�6b��Q���c%�0�b�3��=+�x;`���p�%���cch��겦<)�	�w�%u���^SWr���m�<M|id�~F��������f[D�g<�ĪK^��ܿ]��Y�� �L�K�Q$�f?ߋ��@��w��dث�ǜ����l�BC��x
��i
R�A��<L觾T�p��wRE���nz��%]�Y�w
�
���b71Ik�!1��k�Ѽ{�m�B���'z�H��c�J�����^�̑e���G�#��������������1�r����|�D��$٣fA���:���Y|IX'�ƟJ�qb�D������ݕgӍ����L,*��C��Se������[� �Z�c~��Z�E�J�����b�!�0�PE��֗��q��9h���,����#��W�:7���ʀ����aZ�&�9�޴����]�$�rp��H
d��
���h��h�%ƽk�HCJ[�[��	ouϯD&5S�.(^�J౻�YZ��?yi~�r�������J��^sȴyLk	�#�Y�d�+���t�3��> -v��^]P6m~z?{^+�K�]���"O�r���>�(d�o*q���^�X�}sn�K_@e�P�k~2AqZ7�Y�ҵ+g�!�xѩ\
�k_rd����`�qIҬ�5��/譐��=?�t�x'�,4�k
b���&���(�S��c�zP�̈�_&ŷ(�
,�n9Bo{�	�q�;�)�%�R-���Ð[�ͣS�=�Z9U7x��@���
h�qP�o�t9p��NJOAK���6U;�l�,"{�ܶY�N�AB%G����F%To���8�|��wI���F�t8Y<��� ��k�M�H7�/�*!�#������2}h�%b��&b_r�`UXA,��*�z@>�bpL��"�=�N��{��Mnv��<[��X7}�u����	F��?��N�v�F����(1��D�Fdܢo^�����H?�&���4ٶf9�/uV@��=�������z�\�	�=�bg���TK�&ޙ/��)HS(���OSÁ��m�7�;ýӵ��Ml�^��4h�QU�w�h��)����Y��W�3kOQB�N�9}�~#��M^Y�;͟�Lemˡ�� ��(QDi፞m�ǔoO�������%�+����Sw�epG���FM�@M��ܙ��,�.*5p��]]�[��O{"s��;
T8��lt4��h\!��2�h�i��%>��ax����$J��W����:8�[����s�>
u���Vij���祿C@2��&7��ߖ*������.}n'o�2���]��y�]׈�Px�e!JPU_���'d�3���꓋�ʏ��t��M�-�B>�+ؕ4w.��F'f�$NP�>��nI���p�$��-�6q)ԙ�$'�Wz�ݓ3��sx{t`�P&�+�ע��.�%$D�V�{��)����\�_~7��������
0���c��pNe�G�
��\Ce���I�8���7ݧ��X�HK'�ѽa��c�q��x۝${k�� M+]�A�������_<j�s�z�Q��.1fIQ�1�V���X ))�Z�Ʉ�*�Ql��JT�Tb%N��*6���o��+��J��Ψ̕~�~�X�S�nb�7Up4�T��@ї0m���'o{6�F#+�G��t]�,���=�z�nnݝlb_,m���zO7�@�u����^�	���ܛA�	�P8*[4W
6F�H��^�'-u����J��	厗�x@�C��9�c�='���¤��v�85`��?4.Eeԏ��SKr)9F��V���9>|`� <'����{1�Q:�б�9Ԁ�N�8� B=3��/o�+�:��� �p�n<1z��>�i���)*^M�ռ��m�|��Et�gC�F��8��('s��:;��ٓ_$۾ ~�m�`�YD�rP��9���[������!�0,�a6�ߜt��¿b�[܆��NLL:{$t��1��Z4�S��л/��۴7�s4~zR�)? ���Ѿ��-�5/��}��H�A�s�ГsS��&N�i�r�y��%Ytr4�!x\T
/�x�
z�כ���3ޥR_&�9��u�������S�����t-�]߅F�6�nq�>�����D �G'JI�jz��;��3���I^5�G3�ē�BOf��{��LO<��XV��vm��ԛ����º⾝��%v:N�,���L����o�8��Q�l�V�}�bW�L��k3`"!����"�V��)_�cϻP�O�9��S���h�xgK~ɰ�h���T�n��pyZ3lԗ蟘+�Cb��C�(d�LP]J�"J�iߍ�.̏�i�FH}��n8�ʽ��\/<�<�P](_�w={B��(����h~[�9ݢ�s�!?�i�;�	�,��4a�"����m�+�+r`(N��+���r͚I�PR�Y�\���\*ܯ�'%6�3R&�՜ć�)҈�h�R���$��`/����L�ٝh�q�!j�� �x�r�����S������9��-떵��7���buN��BܰM�N���;ɵ��v�2P�듞�/մ)]�	F���W�u�������W#�o*m�nY�ã�Fs�[�r��n��#�`��А��I�]�Ѽ�k��`��ҍF�`�s�M�����Z܊�����n*�$㠹0r�Y'�[�!i�w��.�	�h2=�
h���`���Y�>�y�����=�v�5�����:[����U�N�����3���m�Gf\��*�)I;$�uz̆Œ.$��T㧺�Kf��A���>_�6$2��l$�h_^�v
����%�?GÖ�GI���I?U���ֆ���W�̕2Ƈ�/xf=q�-A�
�_�ys��Ț5j�jni��=�,���b��Z�NFi>���� �\�v�q�*�>0�7�G5չ��N߄)gF}�w�
�����u�@�[�U2�e����r��C�@:hE�!%�e���ϗh�~];B�ˁ����t��K�N�q� ^Nc|�gMs��*{��R7��.�o�9Vc���F�+j�hc��a)`�%y�t�	L�V����t����+ft:dR��� ��))\�BR��Z��L�΍2M9-��Sf�Fr&�����i���3�r8�l21����f������)ܹ~�`e����\bhi�ڒ�U�7g�l�fx�=�E\��2����v�r4�3{,�r���QQ��*��4�eV�W���^r�u,a��$�e[��́H^)I��S`}B�@�N�o`�{��Z�6��@auW 
 !tn^I�Ě�T�mD�mc�"�9vu���oR�uu����a��l�:��]p�'������_df�g^�F:c���i�e�������K7{�b���+ 5(Ȅ&x���i0�{T�&gE�6�]�W�v.tW�]cNV������uf���\JB�'P��h\�9���ObF55��N��t�P5�u�n2��!��~^�٧Zp�:��.��.���(�hBg\��H���"��e�v=����?~����c��o���o<w����k�����>��/ ^C>m&�h1�4&�~�K���d�t��&a8J�)Ab-����������K���vT�.>�웺<�F[*�C��oV�5�7d򼦴=�d����|�w�O�),!�|����f�)�2
��q4�m�����+u�;m̻�ro���uv�^��ق�����F7zʡ��z�2��>���sҞ��] Pg�9P2լ,xwۭL�<���Q���B�|p�\\��R<�܎f�iq�B����S��W�;�;Q9j�7�?� ��ί��x�%.d�"ȯ ���99-�#��V4S���������c�b���u�����Z�h(M�1����L���Pj��q�Oӻ{�����+��Y�W2��F��eP��GT(�e�~윭2rT����ۢ��>�q]3���3���=}�d�;H;�qᘩ
	)H�|ːev��VQ�x���χ�T��p���kN[v�����L~&�|�=��>��䳜Ҷ�=
8�b;4ѡ�|�Jv�Z��9c�`���d�^�����T�3]��&�޾Ֆ�ѱL|����4�>N�%n;j)(����@��Ǆܴzw���,_=���;U}/�n��Cw	���3���G�H|�2��K���t�hWU��b����]�Li:�7�(�ӆO߁NPD�&ѱt��q���iD�c�?�)�y��͡��kl��W]_�%aR���N9K�����ܵJ��[>���*^�J6�)�HQ��0�08�2�tp�����򪢍�}�^� GM<�0,h����s�p�Ղz!��Ef��b� Rw�J�މ�3�7�(�T���5�`;}��Zg����J�Em��\NBv�ҵ&�Xu�!G���ݹ���Zؤ��KpU*��}�^�|~��t~�J�"bo9��5k8����gB5G���<��jju��K���Dk�?฿GJv��>��oì얧��u-�h��������q�ܚ�ˏGV�B�E����)(?z��}�4��ݒ�='s��P�v3��P�d;b��ע�~OɈ�YV��z��;�)C�n��������iG�ǟ�aޜ<��(G3?�0)�g��N�Mտ=a���g�����A'Y��,0���`
��C<*?��?b�z�1�	;��Ҭ���A�b���<�*���H�GgVV��}TkӴ���4#S�b˘d�%�����ya�iK�N�%GQ�Z
����f
L��|�tFx*R]X"s�}�=��wz|Yd�s�Y�r�u�-;��/lҢ��v�!�4_&E���8�K��}��M&7D7č�q�Jߍ�*��h ���Ty��fUh�VI`"�R ��)��-���,����.�A^�ƶ�����U9�
�&���"�K��Q��$K�&a;Q� �I��J��\{Vt8��J�%��( �Ŵ����xU�A�d:�;a���בfg����`������j"��֮��3����fZ�9sd#�?RyR<�Z������Ó.@%o�!æ�v�^_���[�2px�f���]�O>|�WP��{��9���6�^�J�z.N�qy�F�ɚ輔� be������¿]Q��<��+��e�� ǽ���w�E+�I9���������/W`�?s��.�h�l� �3xm�m�+*�%�rL�_ �[� �S�v�Sxw��?�X���۟'!sw� nQD���9���ބ�q JD��㷷�AAv�'����V��G���㵃���#�6D�
�y��_�QD��|�@�k��WZ�s���_'Zh����-�ݣ`%���/j)>�/���)� �m �4ir�=�}3�i�Q��(^����~�rN�d����,�!n��.@Qv���X�<�h�� +�#�@�9�_�]�/���2�@�-��`�c����z��*A�%�R��+U\POjy���W�X!B����P�/�q��L12������$�I׀�bЩL�:8��<Qc��e�����W 3�n%�xYxm�v�� ��=��g��j���n<�a����a*�Z&��Ԫq��X�%>�V
�$�s��'˓�$p�ֺ���8>O���qM�ɝ:�>m�2)����R[�J��z����]9&Ǧ��7<{����4�	9����u߅2���d�t�qW�q�����RĲ��Ѱ�����G������zx�6���D=6�W��vAGo��-�KST��T��":�=����c�w�G�AD!�6@۶ߺ^���� ��Ilǔ��9G���G�ws����|�I  ��[G{_��T�T��"2#e)M�.�@�����C2�qx�4�
 ���)�Bh�a��]��S!�n��Ţ��;��0b}����tx�_HW��a(�i�/��>��d�4�ӥ�Fivc�p��1�aZN�����V]�;S	�̈́��fY̕	����� /�=0�]�Ւ�&��uhk��]��K����:�)�(7�Uj���+2L�2�̵�_��o'��2�:^�;P��Ysy7���+�^��+.ԓ\R�l
>�d�s��WnY.?bӰ���{Xi�7��ժ$ݣy޽E.)�Av�{+[�R\���X	�~����U���,��Oh�`1��oIp�����b�U�ݷ�5G���`l�hS�׍kxb~[Q�+5�`�at`N�]hT��~��<䑢1�o��o�kW�,6�'�����[a�U����j��T,�z��I�T���;�*�K�_�O�G�o���p��[�e3�dǄȝv�i��O����b"����e��Z��]W@!��l�>h����zC�D�;Դ���m��M��Ǟ����x(���<j�	�O~!�#GV�iѸ�\������H�]�Z��=��⩖+��it�~F�X�8���WBM��_#�_��M�~��na�ɱ�PYl���W�oR��߳��-������;O��M�t#��u
ݲ����zw7�.E���1�=k���2-m��uQ��C-�Z:�.xFg��B���Q��w���K��q�0폗��
t�>��f[��Qk��2������sIY�C	��t/� �=^�u��Ga����ǝ����m{w�[�NqC�Ko,��4�/��k޲Ԯ�~-SD�" ��,��%/���՚n�ocAz�Ú��@|��K�,[�l��	ÍJ�O��)��@��m���)#�Fl����'G��g\���ix��+�Dޫ<,\�m��}ux�ʺ�5�I�D���R�Dy#\[7]���q$�D?��������Ij|$�6PO�)Ց��KO#�U]M;	K���}���Uʗ �PNǯ/Ї)Jz��{�|H�̨��I�#K�Ȁ�J�R��׷���$N<�b���z�Xt�*�D;�V0T�<�0�@҅o,�JkV�9@˺��8e����߈�F����cM��n�����F^D3�S��|?ٻ>��z(��~��񬇗������7��4�L}�E>JY�W����t�r��_���ü����H�`:�h�L(c$�� ����J�p�k 5	=)��?�	~�?��K�8-��D�#�ɮo�E�y9�;�f>�f����Q�My�v;?ҥ�jl*�q�)G-�C��|�U�?-�,��(�T�=��R"�^�Z� ��̋	�
���OJ+�r)��	�9����K=֞h�T~�I�7�����R��I|��	٭�e�.m�ˁ�C��Z8����~!$I�+F	tM}����++���
�Y}߲ܣf�q��
T�c�.+j�������]���T�����6W0vg��p��7�^���=�W@НTk�h�=q���1���Aʲ�u������'���_u��.O��Hp�L����>�n;�eN��}L�I�BޣW��&L�j����
�qy��c�kO�Wʡ@b7"�:܉Bh�l澘�j���?~) ��HgOl��R5D��G�t�
M>��(O~b��\>����-J���!��@�	�Lÿ�T��,��3ʗ�^�'�L�� �E��7]�{�[�E�E6 ��Fz�}�����ǫ��O�ɲ��ֽ�u;:��Eg8k�*�W�ڂ@���%����z2u���	��]���6Hb�^��RJ�u�+@���d:�̀"2��$S��0>��ƛ-�
�Жq����	�3!� #Ѱs-�d���7cv�{�g�|�>8un������R�ca���p8|803��V�ǝ�R����?��8��V���VxL��u�\�7Cؽ�F1��p���@W�d��c6Y�p�j��S8_���f�r����rߗn�o����&�/�s�\���p�&蚰z��ؼ"�q 1���=��X�K`̔�OH�O���>_�&������#��&�۴�C�.�QS>^�T��N��$+��
�9�Q�[�}�Cf���*IC��G|#��?�'��t����7o��R=�̕�OX��s�Y�j�ܩ>���)���K_7����n�mN
�^گ*Ḥ;ạ���#�+h��GE;g%�Z��8�0o�����f�U��`�а��m?�w��a{�3��������y�j|�=�>�P#��UR�q�����&��]��`�����n{��+)IIi�e��E8)��Zv�,S�{+�`~��.mN�����{f�M����)�I��w����q����`��X�XE�ʪ�Pjw��$I6�K�3���Ku�9�s��`�}����r�D�<�a�m�����.��bo����K�jC{>�F��dj��ދ���rG���]��g�LC������&F�g&)@ ���?�h��1��y�;� 
aZ���l G�q��Ž�>�W���i��#�1�B�N�e�Yq�,��ݥۨ��Z@�^�_�ߓ
��Յ-���!���0vly#�=��,���/!�&?�F�>�f��7�ǌ��"fl�k�u9-�v{�;�e	!��&ܻ>��Z��ۨ\�O�4��⥽��� �ת�AL��a�ė��p���j��y�)u�zm��dh��^�Q�����Ye�$�>�'	)�������'~?_�J�T��<X��A�7�>)���4��Hi��#/��.�Z �`�B�4Y��a��	��-M��F�{��]t���l/K�/𧘲j�X��)T�>J��������VF����<�`�1�m�>��þ��C�s�{(����7��G���y�fs`�`��gYz��N���4��p�OH�骕Fo,���j|Gq�'�瓫��ξ{n�����5E�i�}?y���=Ǎ܍Se���k��߻��
	�ג��v�v��u����BaV�D�L���B�!�w� Z�H�B݀Nݭ�MCTd�����dɼ2�=�J�"���N{^�AjՕ������~�Q����f���4M=4���г���m����� `[.�A�_<����@��6%����������))6z�H�O�黿'Z���>I���T�<���e\t�'�hv��mj@ԕ��9�l��;�FE")D����,��ھ����y>���
�k����5�l�v����d쵱*�Rݣi@�[$�[Rjc8���"1�.ͼ>�*�Sꅁ6���D�j9�ʸZ��6�Qf�9��	� ��;\}޳~|��Rh�Թ#� Ymz���l�T����������21�ٳ��Ψ�nv2�}v���@2k����������4��-΃�S���oױ�]ˣm��B{ɛ��gJ%����� �VW�[����P��
�K���m�Y�il�"��%#_�����*�u"�@ҙ�H����3=]���8�)�ʬM��������Y�\㌮d�L]G��!�W(,�:��.�4-������]z�ϨGT�`���*p�o5(�uc:|�#gk(��z�PW��4��S�ɮg1��/[�-s��3ک����Q˄q��R�B���_R<Ǫ�rUD���is[v��ʑ���+؃X#0�n����li��_[��wg������nX)�2���V�Ü���!mGiDV��tq���v�-D^W���@�MJUQ�07��.�}�ָq/���u�X~����H[�s�����n�7�96ט���;$���,��뉨���I��^o�hM��ޏYX峽�m�<�ங4�������s�[���s����9���<���} 흓��1��̐a���K�@�8��%�7'P���Ye��1���U"�>�Y_�q.��ɫ+�p�Z�2��RL�Н`��G�>��5�n�`b��b�!>{	��t����x��ޙ�ȟW'�^"k��s���%?։ �P�p�@|���O�����q�Jƾ�l��M�Ӵgg�a�$�_�^j�F���6� ��4&�X/B��	!������p�eg_��XxՓ��M�����W �lt��3�t�_颩�������k`GR��&��}���}$��_4�噃j��!Vm���+W�Ki���xy^�Vi���%j�Q�L���`�����~����0fb�+���I�u�����t�(�Kt{�BS��	��<zH�b�P�>[N�77J��f�L��Av�\|�xY�6�z"�-�M�r*��G֩'�(�Rg���BG'"|l*��D{���)�޷�+�f}�K���+8���`��#J�7[��nխ�FAX���XiOI�B�'��L�e���R�������*���[%�Ԩ���Ut��sh(���Ћl�����S*�1��a�R���ؓ��M�It����I%U1(IY����<	v�L%�����y�!�6]ۮ��Q�f�	��<�D����=YW%6��	=Xb!
wȤ��u���O�r���-�,n���w.��Х������;�t�d)�Ł��� 4Zӓ��Մ�,:�ㆷ(�PX�v�Ra���$�ߺ6eK|t��+��!B������;J@�W�My��/�:���W�$皒<�^!�?�?���#m�5+H��� )�)SN��k�T.:zـ����ҋE$I���:R�H�U֎��W�]��R�;q���d�%O�*�bkQ�>�(�x)�;YbqQ��(���9�k��-�-�����a|%�*�.��`��1?����(��pU�Av����;��\�����G�1دz:d��+3ہSF:���+3������Љ��x�+������h�JKׅ��1��Sq�8�ʝ��h�,���t��A�=ｗ���F�p����m� c铂���_����.KRu�������PP�����wp��'^�_Tbʔ�FmO�(��l��F��g�Ϯ��M��y����VG�-��JW�
z�>c�I�Mg�B�d%.M6�;�����g2N��}�K)+���_���y�=\�f�%R�r�X��-�by:�����j�kµC��^<hq(EK!�w(R\�Kq-�N�<��[qO�"�)A�C �y��������^{�̵�{J”�U�Q�����4�K�S����ǎ��{��4�#!Wׂt&��o5�?�NLx��#��̈́0�@��+K��!Op���4ϥ"�V|��
��{�l����X��<�<+	�6��#@Q7�C��� di��-!�@t]��݇��JcEN����b��c�=:�Ŋ�r	I�g?3y�����z6��bް)C��7����o��X�o��&V�*^$�����j�3���-�"}R�M,_�kx�?���6�)����{)�\�>U.2an�?�KL�l�]�����rОVY;:�OL�;���k�E��a�� 4���kB1B��jG� D8���N��zh/[#��og~�TCԎ���xN�xx���
:�ͫ�h�Ͼ/�
M-�,l����A#�A�A�O��v?'tșwP�d�*���`E�� XD2��]��&�M�2��庽]}�<p�{/���L�����9�)f
���"�Г`!��-KH��@��";Z������H�[�R�������5N}uay�+���X<j3wG��hO�	H����1��:+/0*,L�`�m�1���u���Y�j�1��ET(�i]Q�����
��k����دn�ҹ���鍙����p=m��\���������|�.��K�����5S�O�h�K�Oy��獃���ϷW�3M���n�65[xK�h�ňZ��Y����k'���غ,�^y�2b�o7]FI�'F��Ҽra��՗�l7�O�9��#ӟ2���%vd&�C׾�q�	+ )O�l����IZ��!g�ġ@��Z�����tx��T�:-��k�����̗C3lh�r,U+�Q��Q�����+���2�������c�tm#��
�Ub�Z�i��qⶹϜ�x��9�#A;�^��?k����]�z�D�`t��d�-e&���Ј�� �T�#�	�us$����$S�&CƤ\�8��׼n��\E�j�ᡭy���F���LTB�y%�@9���?f/+���Tש��/|z?|D/i��^^QB���vcJ�rM�zw��?'>�����X��\�̊�6�"F`|��Ru	Dx{Yc�
��ުK�[?�8�O��r#{�e+v��p�n��%@KoI��X�i�]���x�X!��"������O���G�l�8-�T������S�/�׻8Ϥ���==ȖG�o���2n���NkM���2�:������� t`�G�DO35�~ح��ƏwLf�m�nO�:CIo�8$��ީ�ܑ8�{�ECD-�Jcj^)�Ҥe8���P�o֊,����g&����@�4'I�)�ubY�x,$���W�����N��4֎�aI�:�*iA�`��0��N��z[�����������
S�T�����%�Pѽe$h��:��d	性�d�'1	�{_<jˌ-�H��YQ�>	�D�M���]�RT�E��2�V ;q�̚���b7&*7bd�yd�r�R�}ט�� *d�I�έY���JBp��vo��$�;�%|�Z��j��ƈ�ȯdܶ9���TJ��4k�gR�Kd�D�}��2$R.��3)h'|u����H8����������Z1����ٲ-˻q�
{�8�bq������H���vby��(g���DH�T�k�'ui�=�C3eO�����R)��I���$�,��Ԋ @c�����F:���@}|��Q⺾M~�dс�	f�G��t�*ڦkK[%�Wuؔ��B>�Z�c���+�C?ӻ���zM�0�%��^ޟ�m8E�(᝶��*�8bÇ-:�����-K�d�~3x�'aBZy)6��=:'f���,=м�g.��0~��T��8�k?��e�^�	�\����cѣ����7k�q�3��W�{�s)�i�U"4���t��9��-D�Hn�T�+�*�=��G��7Tf��Y�EI�{RL�Ld�vO�k�j��*��i��.:���a4�'�|���YWXSvK>����"������x��(������Ψl��Vf�߉�;���3�l�m	�r	�|Y��;"Y�z�{f�x^�j־����8UoH�O�r�슂:�wh-G@5Ja��fW_��3H���?,HE��L{��=�.��y >��@wf���5�z	�y���#m"�7}���=+��6c�9@;A�A=�kO�A��ʞ^�8+��0����ҕ�{u��B+�QO`����?t�[��������O� ��fN��oI�Z����%��%%��Js�O�ߐl=����`�[����1�_���t���t���teqRF��~UJq)JG�'�Ǌfgݸ��K�36#n0����	�� ��Z5�74~7��*��IN����'�j��)�x��:�EljC�?�78�@��Kr?�/�ٻ`�h�{�S]G�̓Y)��W��$��RF&6R�s�]˘���z�Mc�b�Fw��l��&�弣Vh`~�|^��Y�I\��
��z��� Ȭ	���|��<�Z��u�w�\C��� ����BDc�$�G�󥝼�*�9��Ͳ����Q��΄gV������d���dL�if�Ƿ=�yDz8-����d1F�-ːI�hE�W>`,1Р,�cA�c�[���n��ZXp���qcI,�^l�k#�q׵�~ݧ�X�φ=|��AE�#�9�*��&�bI�~Y���������Xe��e�VtLI@ӈ�䘣�X����ºh2zB? ����B�d8�3j���_QUgo�U���.9����u�u_�ڠ��P��Ŀ�V&���2X;��5�N��<�Gx��;UC=H-x��/��4~�ǸCł�Njq��^�!���wB���H��G��jJӰ7��`��2/Â'�hZx[Uh"`�����@`�E�[į����P�ǋ��	4|�t�'�n��Lߨc⠰��~�;��M���~s3����K	��j	h�[6Ȟ%i�����}�FB]Qx.�_�陋��Q��i�������8��6aQ:_�^(��`�\ް}��ܮQ���Bx�0F께��{�&��[�8��(t����*OX�z��I_��&I��3�U���I�=�J�M0�� ƃ/$��`�M�A�<�!���l��0�0�\Qu@�`��H��zs��_$ז�����Ҩ��D��
���%�]�L�X�i0��O�S�c}�$���O͏L.�Y�>�1Ѻ�����8TB�K$�}m3�����F�����>M4�:��u�Ŝ�����WǇf�?@2/ `�G���uc���ֺQ�X�j�ݿnO�b�$��=��}��� Y(7I��Hr�=l�M��I�|�*���&ak`�/ٖ[����lOWԁ@;*���� Yݘ�L��3+.��5�pK����:��!��5��!EI�Y)�Y�s��Xo/n�7o����8(��G�˛5�i}���Pa>�z��($��/�a�!mm��緷�dq>����8$r��̶��^�sj���UC�H�B�&�j{=���F.�8�R��ݿ���_��֫/�-���`��|3f���7O\�N�`�x��ruX�g�B���>�����SZg߼O�4	;C����K?���|a���6���6�9�>��l�A�I{uV�xsw.����ڏ��^��K�Rڽ��3���/�a��o����b���K�3�ְsL��"'�Kc��k�v>�3��,c.�i��6�J̟rn^��4���R���Y�����Z�iYp�Pi��7��k�T?����+�,^��~���s|PF-�D	J��L�	v�(����I:(�Hu;4�QR�y/���;r(��@��W;'�+�D�?K,"�u�q�����\��2�|��l,I���$��<k�"��Cu�kLy�A9�n&���Q��4��2�@��Ȱ�������,�Xٳ��c�_����N��s�+)2=�m�le���`IL.¾�*�ves���5+k�'�Ϣ�Y���j�ɸ'����}�Q�k���,8��� PM��@~Q�o�]��l�#���-D�k����߫N E��(Y=(�1��]�c�S��'6z>;ۿ���=�>θ!��fA��MY9�p���Ĩ��︫|�	&!��o���`E&̛؟�[�r��A&8*����=�Wf?J72�%�Ԛf~�ҵ�e�>j�\Z���lt��_t.��	߯��-�%A4��?�ÿ�$�4+�pa�|�#�v F�h�hJ�D��|R���T!���V��s����0�h*�3���j�.n3�j)��˜|�ݟ��G��c�U&-r�XJ4G]�����5�wXGb��D����u�?���w�s�3V+G+y/�d Lb�</$�+C�YC����-��4����@��AayNf����=+�0Ώg��q�3ܳK/ �2�����L���
�E���Ӥ��q���j���狏 ���;k�]iN�g�)F��\�F�(WǢO�{���i�������h�x5������5���,����ӝB�36w��f,[{���N�:�@�v|���(9��R�\��%;PM��ѫ���߱�f�K�(]�m��6�h�#~$P�M�[DB&�py�ث����T)�Ź�833���&.Fi�I�R0�l����f�P4� P�����p[&����Џy:��Ŭ����K��n�8r��U_���;LmYh��GXr:Z�$H���Yu��[��|o+���Z�0��z�X���� �V�@�:�w��z�X��?�0�=��w��5|�0U<xq�Q��
���4��Y���;Z�F{ȜZ�����A�Qc�%z�q�%if7��pZv���Z�4�8`�^p/��w�J�L�Q9�s��P����������ә�nEiN�r�,v���<�]�����?���^���[�s���Z�	s��Re?:��?�����D4�H�6Z��9�˦���R�	�G�ͽ����Sףڅ���x��C���0�>jeb�R%�MKL+��"'��<cŰ�a���k4��#�(ŵ��L#�#��M_܆"S8.a)��!������'c\Nd�����<��1�8\�\��#��a{@�c��^��͇n����h�Zg�p�i��<�_o�J����y�y���>;�p���r�_� 4��$�.��D��&N*�~W�c`1��ݵ�&��ք�<YcQb�p�j�hN����ZTq�?U�׹�Ršo����V�m���k�~@>8�dؐ=���]ΚHj��̍*-Nrl"I�����Om=%��0����n��D���<@.��E�`}%kg���~7L���ya}�L�DK�[��M/>x�Y=.'�]n�O��jґ�vA.�����|J�`����\Vv�	�#8�d��H�N��->1s���Bo���d�A�'������XŚT�q&2�(�(���6(��U��b}0Q��MĘn�>�C���S���r��6	|�!�K�������p��ȋ��,P]8Ld��w��"��=X���s�r�V�Rp��'b*Xpd��4�B6l� 0@�_]R�𩪫?~�91��a���k��W����|��;��[I�r�Fy������E�~�Z�K2
�
�!�a��r����Y���wv���]	�d��]Ǽ�{u��U	ïS�k�Wi����Z���:E_ ����N������0��2� 9r���K��Yb�/!�ƪ�^�ݓJ��LIM������\��z[��Y$���.���|��`����x�6�w$ȡ����$o/f
ՌK���|����W�/�á�%vU�%�0�њ#���!���+W���G-�?�S,���4���.��)����j�ʽ�E�U����G�N{cT�4� ܌�<N6��t�]s4��﵅�c��Ż�m���tS�F�v@{�]}���%Y^��|;��Vi`I�B��S,�I4��!��{���_�%��_��(��P�Ǥ�m��߳g-��~�݂5!,���)v�w��8׶�'0�$׳%Ѡ�=Bе�R�N�iZ��5�*L�!�F�X�AO��d&j��������8�rtV��������4��JǠ����O���M�5SIC�<�NFP*E��*��a#mR`�F��fm�&�0zw&��6c�f���2�������P�b%���2{QS�>�oL=��o���ų�-DoA���A��ug��W��왅-�=cj��;�?��Q��UZt7����$��f85�_ !���c�\�Wa��^�yv��yp)�A���V|At��˳m��e�;v��G�r��W�]��Z�*J�C�'U��:�F��qa���\���<���[���b�Ɣ�=�g������Q��w��Xh�tM&��[M ��0�- ����3��H�'�u��^��� ���4>���	5vS<\�)zr�鈮x�#D�;T�Qo����bn�r�DM��@������t�|�����S����Xp7����A-5/bXv�i$�ޏ��;�2Ba	�֧����*��j'�����+���n�-�>@%�� �;@F��� +���l#���'ai6t��ҏV�� 7q)m�7�~�׶e� oy2{�q%�<O�n`~�=�!�rd��g)�3")��~O��d����8�Ȧpr|�rU�;$}���@cv�	?�i���Fk�_�I|J><��)�"I������5�z/����j��W�I��ɔ��J���k��C�7���NxM�I�!2
Z�)��~�PPb	�a/UJ�_���������o��� <���Z�4a=݅���D<~��I������~��9[��C��(j��m?J� x�0Y0�E���OJD��:�5�*����k���s歹t���T^�Kya��_�4f�~lb�:��0#�[�����Q��l��J�^v֝��4�N���Ded�é|�py{�t���^}�DIܤ�O��t��u�<~���^�G������7�����{'�8D��r�_ ��m����!����Ϝ��9|�]�>6�e�>p���?�q�
�#k(�>����}5�Z�@�ӷa%,�.�b�(�E�P���@x@���֬��^z��m懞���:�G�?G�A�TT��B��Xb�x�} 1��'>��V�	��Bv�n�b��/�vc����&���&c��� ''���
�P��Үi�ҧ	,tE�L��1ѵ�d	���ݥB5��r+n��� �*�|�!ѽr}��]u��������4z�V�L
�	ڌ�R5����ytQ`�R��N'��3a�-�\s����VcV�c���g���(��t��v�>��s�QPJ� �	����ٞ��x[r���o��&XA�� ������(��]��17M.�١�� ��ߟs�=}Nj۳.t}t�Q�h����*�*��UId#L���]����]�ծW��#<��M̖�t\)�| �|�"�IJ1{(����y�n���0�9� HO���dWP��ֳȝ�^fY
�� �^��A���4�o�Ѿ�E�ۓ'X��������]��γ�E:���e�q\�'*c���4�D��b`R�Y0����Q��.K�o�mQLE�M;���C�Q�Lh*������h=�7�����n�
�%淒'�R����y�}�6���~�|��������<OB>?��p 2��v�/J�:a�ĚO�hjk�,\RBB!TJF)9W���D�Q���胂>��ߡ�����W��[���Ȓ��n���P��=�=�+��=7����T�"k�L�3v��W?��AEX�;��.x�V|������^ݼ+#��#"����E�R(��fxƔ�m�Ӗ�Q�c~�^�� �YT���j�#g$v"�a���sڃ��σy����_]�O�[���h�NҊ=�v��r�Y2�6��q���)�ᛳ�wnQ�УQ�&�y�A�s��
Q�$G�3p�y�~������s|$����g�?\l�.Q�ל�c2&�^p,*YC�8�i�Q���Yq��+ox{�G̷H��|o���Ӥ�$���^�e*����N�	lՃ�w�����@0�����~#ͻ
L�!ěuR�
��z�q	-���n7��8�����`+�������|��{��I�$�6�xRz�*���O=�i�>���c�J˂d�E?cc��v;J��v���Ș�9G�����}���u1B���k;��T�ٝ�;��I�P)j��܎�B��~5�^R,��~�S���U�`��Ȱ��д�6��m2u�OTdj�"��:����~^���),	\k���D��f�#h;��	������9��R�$1����G�p��"����c�o�,�������0�9�����{XZ<<�!�	`w����X��A.�ZKf�sC����~�QOPZ�?-�0Q�'�b�pc"$X��6��Mx�1�&~WJ�g�	�
�/
Qsꪔ�m%��
�BS(�K�ޢ�#*\H�)���a
�\�*o�����/�p��s��I���W<���]��YmQ�N��m��4Hb��ʣ�f8V&�OI��2�݇i<S�f���9 NJ0�"<q�-��ۺ KV&���LV:QO��L�{�*�ړ5ʯ��'Юx\_�0-�n�)m��
�\і�)�ݖ���%֌Q}��X�W��`�|1�Z��XboWK�C��s���FMW}2�{���s�'R�o�p>p�|D���t�P�g�#<	�:�0��x{|9��̔�>�V��^���l7~ 7��#�)����fk���mlE-�U��k^ k��E��;���Q���wd��xL"�/ ]?�R��h����2�&axO�\-
y�o��XvX�-
���7��F^[BF#�����ɡ�.��1an�S)��՝��Q�u��=��������|E:c>� �t�r��u�0�#�zOZ��G�Mq��ؕ�k��t������eV)�|�{�֭s���ks�>�r�b��T3P��ϧ�Ω���'_�3~�dk��q�O������=ND�-~�
�λ^�(�S5���F��j@s���Ѳ���cy������>1� Zw*@�?��۪���5�cf���$ɭ��<&�6�2��+T8x���sKb�8�oh��p�Rt�x����Y��d.�t����4n����h������H����5��{%Tɔ��(Ӝ��p��_�m93�p/)n���V�ko'�(\��(��g������:�ܙ;,&�׃>��f��`f!:_����+�%�F!ŭ��y��ƪ����^d�K���ER�z�(Q���N��gI��'#D���@�M����!m8%t*�q�=�"6����Ī�O�`j7!����}�SWz?t���/�l+��耗�ܰCj���2װ|�ȿl�[��ึ���#���s�y��ԜЮ��� LJ0�$q5[}w�����gE��Ob�;`��֗OU;�a��U���K�X a�\@|EmXdS���P�$����
��79#�7�Tߪoo����7�QW>~�7~ZXZ)dS5N$���kg����a��NN���,�q�o�q<O�1�?[})�}x�Nܝ��=�R.�u��Oܛ�Mg���z�	�^�;2��Vy�r���{��|ҩ�-���#Ǘd�)��,���Lج��'o��p����|Ł
<"�Y�������vP!&m�x���x�;	�V`�$;�N��]��X�o"N@"8��x~����t�b��}8����NZ�*g�1Oyz0
��R��v�bJ���:�\eAa<P�W�q�M����'���W1Q�8%�˔��ُ�^ �?]�V��<���{c���>��Ii�y.ޱz.�F���M>�TK���䧩�­[f���{ٌU_�����S��ϛ�mg����o~�
�h'8(n���h�~��JDaS��t� e1dN�A�\ #m?k�픗�[�k�cf�(��қi?���&+���44��P��5�=k^P��@k[y���i�_�k�fv��|@�*{��]uʯ�4��c�il!��X��ު㗖�r�_<T����n~��<�q�?�LG�Ӓ��	�V�6EӸ	���q�e)�} ���Q��r��t;�&�?��mV�U�M�1be��74�{L���.�M:��u:9ɲ6E�d�,~"}�A��]AG�)���υ���h���v��1��x��؏�c���������M��)������~<2L�/��{W4*�[>���b��
0���e���*���H#�CJٷ�.$s�Gqs�2���,���;'�TG�c��'�~�k5��S��ևC�3��s_�ZVs��}�dk^3��9:o���%�S���-�w�t�=�2=��?:�1��[U}O� C�/^M�Pff�+=��H�e:�u�Np��Q��l@_T�nm/O��g��g'�!��bX�;��x�Xq0����P�fTqVH�EƦ�(m�@�i�=~K4ヨ�&����m7�=L�����B��k?�JI�a�8����Bؤ�J$�w��ʾ�I�`��'��E͡�@��c���A=LjB�~���e R��d˜vR������1ĉ{�+L����1�N��ny�ڒw�r*��l䗒d%�+��@�9P�;wZ��B�5�}���'�fB��Pv)�6�u���h@w��C��SOk���Y^�R�c�7uKo��̢([���!լ���V~�2� �$nY\g*�\^�#�-�w�D(W!�r�Y�u��rN �@	5*O�x2���cg���e,v��=�W���Kiiz.;u�"YW��� N����88�'j�o6����i�ݦ����*<GL*<������ �#�v�e3}��G�����CRm�L���L��9l�=Xi���m�灉[�%�ן�J�1���FQPmF�5C�n�P���T���B����%=�_B�
�O����^G���?��@�����!�u�ȫ�c]i��J��g�v���@�� έ��G�k ǳ�~��?w\��z��bY�J�tr�|B����z�y�~\��ć�,_�q�l�y�]O�L���0~� ��C��yDO��x�@�q|���&���gױ�a���Oy6kzR(���qH,V��d��`�^C��]w�L?�骢���Z"of���G5Q18>�w���u9��ڷշ���yd�1����BXua�v�D��ӄ4g�Q�h���y�{��%�J�I)�7{�m�e��;͈�>�\���8�Cz����8x�Κd���2�oC�f�߇�"��fku͚�p���P�cR.o��W�i��.~�+��>��;S��gG%�"��b��vbx[�_�h��\�'!�H�	��������ߛ�D��nLT`�.����{��tӼ$-�@�4_�M�XĆ}M�.���ڱ�����y��|_-���ߢ�¤OʷBR��,�ͻ�L�5����u���u������{�a���r9הB~ڜU��hMU��3	^����ķ?����كZ�]�5�g���	���Q��o�����I$�	cey�"�@�A�6��������*�PKX>G�j�Ck�ah�?^������I��|������V�
i�Z�[��m�P��F�jė�.o��.3w���$�,������c7�њL]��񈘭U���B���;(�j �W���w
�b����J$8Fs����,@�����g{�Q�\�
Wf'j���P����D���#��P�̾#Pc�EV<��CC9�e�>��j�N�����ʆ��V+}��Xm�t��ɯՉ�.��
�0�F�����C��̱��n ���e
-����Z�CWǎ�{���-���ߥ��䫑�cp�7|�<Zr��ƌ�(�~f�G��ZV|�C���)��ǗU+�AOm1߹�HG�
�piӏ߉'�{_�����/%���K�rmW��N����ٞ�-/���y�+x���_O�F[r��!�0hPP�����MLb!��=q�rgb�3������C����3!�Ǆ���/5���Rh�A�к�7�DDR4��qtgӫQP���E���Ԉڇ����_��g>�)L�c6���t:��G�/*��}���EKb��)`NS����x���]����固�Mk� ���u=.���sD:���]�98��� V�,��r�6r\���Q��r�1�Pr�puo����m8̡;V���w����up����X���y��_[`�"%G��+xg���%�߾�e�*�^0��<��l� �b����~���׏ipGeQꅪY��̒��\!y� �m��hj(T��O�嬜�[0�1���1�x���KO�/�__~&���:�*���l48� ���j����0bu����_l|㤡��\���"!�&:u�Oy6$��"b����+�]0�{3Ҿl�1��4J�V~� y�!l�/C�N�35����Xl��6�u�&
8�{�5J|���_�6)��|�Y�h��}t���t6v�H</��$��^mjGp]ZD)�.�x�`��kRpmL���@��?�^OL�v����Ӎ��h���06G��a!&�b���|��S��k˓Y�z(���`��gs����,'�r0qV���t�y��HL�g`�l/�du%!�}dy�0����y������=r]���_cG�6{�{����VPi�-Oi-��{����	c{f��Fx�6]m�,В@X������6{�Z��g���x�?�*���:s[�·�Ӛ����G����Ƀ.O?Z�#�ٓ2X���ݶ�.��*���ޘ��Iѝ���,�����W`b�����?��;�|C�)�dv
���Bk��U�e"��!~V���Y���l4q�&�<1�򳬂�;�%�>;�_Q̇�Ks�u���pcTn&n�[�	(6��M����͖�RL7����/��VaQ�*r,^���>�AV��F����W������j)�<i��4x����dD:SP,(X�&V�BQ��V�^j�nm �2�'�4���՗a\�`��Qz�w��FbM^[�H?}����}�=��Bؤ�0���� :HI?��D^��>���p#G��]��c�.�ԗ�k��J�G{�N�8��WQG�,������lJ-������.7ݟ���?� j�+��Kյ�scO��u��b��Aj9�#3�ԥZo��A~No������2�E�x9����R�J��{^ ���#RlF�j~3�QѨ�~��`�Ͱ� �g[q(��/ՄՍ��V�1.�r�뛵Iw�w)�2�Lb�NCrɯд�K �wi��3wS��wF�W��*�&4 ��/}���{[:5Y�l4T�R�4*}4����B��e�A��ԝ���4?h�}$��o~�/�X1T��`C%�B,�h���+a�B�?Vb�2	�fo�ܚAZ��;�l-���>�PJG��Gw<�+���C��^C�ݧ��x& �"�0����ʣ�7���H-�	��ST��^�����?�a>6��m�i�n}Lk�r�|Ǣzt�S�eߍ��S&0^Ojf�o) ̫+#�41#�}6�͎k_Cp'F���W �?�+]��U�J��tIu0Q�Mk�!��!�˃�|�e<�y�\����/�6-ִ���>���r�8��2��_s+ժh�������BF�bؽ:�Y�s�/m��>J�'�ݫ=<*�>Z�"�-�kw.*%הוB���U�j�V.13��
���.1n.;ٜAh1��ؿ X�pخ���x,����c�:@
�WY�� ��l5��u+G�9�+��N>�<�:F�O�R�rU�S�+�!���@���˂�ʼ����L�J[ξ�6��Y�G�ˑ��/#�ta:`�VP��G9��w����ݰ��L%v�:0e��E�S���$��4JIj�ގ��ɏ̤��͐�l5��KL���X�cq���L&�֫~��q:&��MV0PB��Sj浛��[Z���OL�v����i���Z�yZ��`��W"���S���~�L���`uK�v�A��ػI�0�vvW�Ģ���A��t�ͦ�@W&�VSμ1l)�ĕ%�1c8�нW�����rU~���:�F ��/G���6r�D<��IA-��|7���z>S�H[8W�(��5���Ԙ+P��1==ڷJ�?�,�<���}�W�f�f��yox�o����@��7�˘7HW/���N�����o�.fH�eV�юO���o�i3�t��vV5�w#p
I�����]��I�}�r�dV2-�U͡C�?���Գ�o�%T#�ˁ��c݀c�o�O���~�4�K8�#�&D5���{l�6��Y��Z&����W�������&m�C�	�"U�4��b�h��j]��v)�D�n��ޓ7�������u�I
������E�к�F_�WR��x��B��%�hDR�@�I683��#j�"����.�8�?�)�c��W�#���nxHHYu)��V�����=@#P�nMh&oN ��mCͱ-�
�d�����ee<��<z녞�H�',!-��O�5̔�&���~4���K@��
7ek��?�K��1z�>�R�Q��,E��UV0�}]KeC�/��&��i�vm�Jg�Q�E�6�9�7\���˼���|�c�LډX�v�57���Ƕy�_�2����
����.�_�|��S���w/�V(�!:�|9���m�m��L�㌵a:�:D�@��Oi�]k�����u��D��'�dw�o��=
�ً�*3sE�{{Y�7b@���t����9�^�H��5<�F�E,��~0����r�3����^��t_wu�ÈM0��]�T��PG�@��gr��&�o6��[N%��w��_�U׻���Dn�����L�9�\L�hs��F.Da�]
�2%+A��%ڹ�Q��7�T�;)0���E�s��� ����#]��)�������K"���
sIw��Z��!h�`�KZ"%6�b � ����b���>��G@*���/2����l�NM%Y̹����@EÍf]k1̩sDp��0�Z���/�wt�F���?�����[�߼nu����!v�V�E�"G>��ĢH���w#}*���ݩ�?�(��[S��{A��}u��cި_�9}��$�*�~1��H���@fK�l*M�/�˺��.R������$�+�&@;��WǑi��Ps�4;)�}���ڽ����:ʩ��O|����Cu�;��gwf�1"Ed��@����O7EN��1�J��� ���D2��Th�S�A��CM�2r��W���i��7~�NR��C��2j��5Th�xd��\���8�o�C���1N�VQ�A2A�cq�|���L�� ��S� � �}sA�g "����GQ�ҁ�yZ�ls�J��Y�� HJGue��dX�D�7��Y�e��o��&�VL�I*G��&�QO+�<I�mx����fr����%�A��f���hI�z�!e�s=p��LۏN3�=�&"˜��j;s�d��赵�'Ϊ3t�h���>��=���&|0*=��R�2����I�̏�k.%�D���i�(��U�(4�:f����� n���U�����m�p���WӜ_vË�"���ԳB)�ǜ2O�P�Gö'�K��W�@�9d��!�dь�Ν[�����ϩ����>�}�~uR��T�y�?����#Z�Y�2=<�]�n
˲U��R�?�Y{4KP>!�]/�Z������:�q����bgQ���)o����������[?�e�p������É� ������xl�}�d	��2�׬I�?=�M�գF���L��p��R�S-<��*��`KV�O��~	4�����	?P��S9�)[w�斳�[�{�1��X(9'�>����	[� ��%k{9�����2���t��;ß�����-`~�1`͕^BZf/��t�y��v9����M�Z����,�uc�ڵ	��Y��G�f�M���B�.�����rDڜ?�,�L7@�h%�aINu���
����X���\�y�uzl�d˽�^{��g��B�g����Viu���=F��;�Ӊ��=��c�8˕:gk���1Q{
��B�*l�D����yK{7�jo�SQ1UnZt`�x�&T6�5�H�0���ю�i/g��;˾(��/� H��t�4���Jw�t#�ұ��tw7H�ҹtww�r�{���<;��̙���|Ǹ��OY&[ʦg��kyU�lZ��g'��zoc"�5�h��e�&$F��1GXsD��ػ�^�8�!�G ��-.�[��Ej�?�y�	
K�PVQr8��F|o�f�Wo���oʆ� R�_e<V�OO��Q!�pyg���-����X�Qdt��O�V�^����;/���_k���M�)�;����x�;M�N"yk����.��%*��z ��
���<�°v�����I��6 �,�����Ѩ���q�yP����N��k�2����.m`��j�~?W��[�}qp�f�Y�ug����f�ใ�R����[[���ʳ X��+K먓��Jw�[޾b��ʕ¬,����0M�b,�S5�:��Fj᯸?�_�O:Q8^��޻�Izp����3%�@��&!	�G�P�`��Y�V�ֲ!�h��코# K���p^^vkN��U���;�06J���~$BO�-]GN����{eqߍy���S�C5h�u�;���;A�z��/��xqb�%�#a�z^����H�Q��Ύ��� �9�w���b�)��FHˎ��Zf��X�š�����$S��̚�~19�uQ������^a�/ir) p>n�<���M�����ﶤ�r�Y�[q(o�D�X��P���N���J�ܴ�]�µ/��fO6��՞��|ؙ;\Gw}-l�w�]�.�i���)�<4b����4���(���G��b��J#�1�KJ�݃tU�-*I#,��k��>F��haX��>r��f��EZ�FԱ��t$�S}E^�\\z�+�Z���/�f��{Ԑ���N��5P�wz��(~����0^gW޹P�KH;Ձ��Q�����n=n8�mE7�L�35D�3�N�����@����,e��ɤ�lc�씘rqy�"��_JX�3��򭈛�\$m,b:^� 炓�ї']5�?iY������t.�晛GZB}�hƙ���m�"s𔌸��0�p_���.�,�3�V�A�g%VcҚx۱��=�L-��AE�^H��\@D��\P�t:���d�z3 `��Ѫ�^B_98��c�E)��OK1O�d���1@�z="s�u����B;�We��[1���/�I*۲�R#�g�I&��zXE�B�$��P����\)Z�<U�c�jVEt\C���,'���nh@V�;����ucJlx�E��rl.��ܠP��~�i�ʰ�W*���L9H�P��$,kEV�oS]�)�2�L�0�$+��ԃ� .K���(KWG�xp�f��u��Vk}�80�y�m�<��c��9�W}��6�:)ȼ����S��E2#F���TQH�|��V�9�,��ř�����A�#��b��>[�ʜ�{��T���Z4g���Q-��g�F��:(��?7��n,~\��UHM2>�(oo���E4����C��kZ��)�l1�k��&�؍�/`OS�Vf�M�)D5�ϲ�7vPޒ�?<8]Έ��'��|�m!)`r���$��[�(��mt����\x�w߭�ݢ��DA�&�bS�MV�i0I<�C�����oT߯�_�y̿nc0=�"-�᧝.;���Z�������boEW�����^�3�����k�۲Ѯ�z��i�S��1�*S�ou�p�0�R:M��K�4�d�S=E���Q9N��y��N�����\2L���aů�
�P���X�X����Ȥcy'��ڎ�{T��h	\x��0��jⴭJm4dX��=�#��`�ZOgcw25'[���+�� ���`�d��Tפ8#E�5���c�#�Z���y�)�T��r�y���XZ(e�	��oX{�_2d��l�Tܙ	r�����-��_+F}^Z�8�Z@6���w�0�}?Ga�!hp�asFyi�����׉Ͻg/��T҉I���ј�bԁ���32�`�x6�T��E�v}�U���tb�(�ȑF�+�v�5���~��]� �p�2�u�a$�$HF�=7���%��r�[|o+��kv�9�� D'��q�P��E�Ϻ��B�?WSy����"牏��-���ㇽ;��z#JGٳ�4�5���\��D��(��;����O���+W�6v�?0�3�~�t��J� �k�p״�LA�����;�$ӓ_$�l܃����Dx�s�KH2���2f�*�|Z���$�x�U{��r?�pKщJ�I����Z�	���:D��'3<�w\}{J�d�ba�k����6��*m�E�I�ǀ-9��v�����)@�0h�����g��/�"���X3?�ؐ�]���܆�}Ϙq��������hG\��"~�.c!�"X�_���/���*;1���K��R����R��Y�Oi�p\&q��$�:s�6���;��̈́>��_�r�[��-FGSQAT��)�ⷌ0�,�W��EjUt+U�>u�M6�t_��
�lG�����4�v5۹}ȱT�����ݖP��s�(|fr�Jx����>��5m�����}1��Q2v=`yp;���2�n?��e߬؍<��{��ܔ=��W[�O{�Ɨo��'a�g�lkf��a�f�Z��Ar`R��y=�\�Ȏ+Z�Z������u�U�R2����J-�󾍷�N�xK����7q�����Cq�\z��D�%��'����I�����A5���� �4��^�"�U�A(/�@N]�����Q��e�H�Dbc3M�獤^�CM���9rJ�25JRO�pI:����ub�Z�b��$s'�G^��Pω;�˵�/(�U�����.��ŕ^KRjZ
=N�0Z:�L�����J��D~��,�"����W�r(e�!���ۡ��R}�Wt�\X�-j9�0�T���uh��.�#^4|&��w��|��2%��}��r�:?j�(۰4#-,-���YE�d�ɬv�-�A��|������z�v���Ja�=�`-�;,�<���Z<(���fXIxKttѷ
�p-��Kz�����:"d�!��F�s��vW��t�<��अۛ��{ں��_�d�f��$J��Ӑ؞����`�������s*�+ R?�
@��\�U*'�p�����!�'�&*��'N�����#� ��J��7qu�R��+��{r�@�M�,鎼~�6��:�"�0��0k��6�=aC&�G�Q���4^���-�&�����F�E�	�Y�'���pz������]O�$. �������J$'�]����2�x�;TA*�ѬvW�@o�R4#f�X�b���Oo]"7�nn�~�F��C�ۆ7�d���c|As[�6C�"����T�w�Z������"�$w�3��H=�^�Qc�����V��l;��]������p��ڳS��i#jchX)�[�2�;�%����3[��(t�3��v���+@�v	^�ÓDџ�H�U�Q������9[�����B��S����_�^i��
(�^H�Cf��c�أ<�	�l�[w�dl0�5>ܦ,��;�ާ:\9^n����TI�ہW�:xp
��o!����S���Jlw�޼�+��$u�D��w�c}�C$(��t5_Ugk�V#SȤ�lR6`���|'-�9�Q��5,�߸,'�_�hգw��[t+�lr4���HmQF\�Ik�f{Z#�;�,�ҽ]1^aJ�n7�ۘ��&�-8r�xd�P8Ob��O�����[(W�M�)�'֒�+����0Ʀ�&k��Z������l"(���,'�ܒ��Ƥb�R�,dpF��(�-75���v�E����K�T�8�+ )W�#�u��n+�]f�℺C�s��zj��iI��m��Y"������C�n����>�p����%��R����U��e��L#�P~�XG L�88�P��y-R��4��>c�M��ӓe�8�X�hk��g�K�ϯ���Y��^Ҭ����@0���^;�a�'�Hk����H�tL/���(ݶ��[�3�����/ �'����C�<�P���cD��H���a�(P
���:�-߈�[��(�ru!�R��_� J�ͷ�Sr��!��(C�p��C���g	i�`�e�;�9r���tb������DoƲ@9�H�Ě� ::��H�-{S�5Qq�yE���������9��	� +Ǖ���Q�ƴ�t��f��A^���g�d���7w$/rauT��a�?����m�l��H2�ox��5����e:v��/R9�f��^l�[��IT��+��x�<������u��w���F���Q�h(�<~�:���u������u,��L�S�o���-���u��Ek���3�\r��U�:{.�Ȣi��h9φ��,�Ȍ<<ז��;{�_��V�nI�Ho�~�.��g�ᝡ+ҭ�����Q�����z�#>�z_�2|H��ӏY	�JGY�	l�� |�N�
��k��s��#��綝�uY.���9`�J��(�MT����"B�Ҭ�C1��_�4��S��*�#GU\�L���0�U~O>ο�Q{jK3��	^�͈����5p��+���e��8�:�������=��O�i>��M��aB��<%Xl�@�s\�����@֌;�XΒA{*Y��C[Cb���@P�ZI�SuO�j��V�IQ.P�t?����"f nx������E&�5�������>�mٕ(��G�l!Q�����ބ��nQ˒��
}�B���OXj�4����iO�r�>���!�C��hOz߫DL�\t�P!���t���Kc0o�Z
_�P�K|��mM)T�<*��S�9UDlG�v�OAHְ�
<W�����r�Τ��
!L|�`C�3v���7�D�e�/�0�[���$A%���j���ͳ3�6K��[%י��C�����f^>�:?&�.9e"��v��N����n��R-'����S�\���/���+�FQW.����?���K��mJ�T��]Ji�$W�?�[mco_*6uxH}i��Ⱦ�d�ǃE�۵�1�vn��㠰����##���`5*��Cv�Xc�{�:hq	۳ݛd�VO�&��y���A����QiS|��JP��+V�����-V�l1/��$~�m$��+�g��X���AV�S�`|��*>O�\'6En��7�YM[����1���m��/T��N��Q������z¨;LL���`K�no)��(��
�EAЃ�|cW��"�z奒�S#
��'a�ا�hMz�3=h\Y�W��Z�l.1Ğ��dX�f��O��u���T���|&`�z�W@���o��#�dlpA��ۚ�������J[���5��@M�@E;�.�@J�Q������`��J�JV�����s�HfM���="�~�L�B\KJ
�OHF������	F-��|@<͔ڣo��%h;�{�XѾ�����N��Xz�7)6��$�9�-�ou/��(#�����4��7����+I���J����Yf	&]ԡ(���?p�����16o���^�s�8�h����3�x����7b��T�|tvt�XY����"�a��>Aw�I�t,U" ��+��X���B�Ի�Y���d!*����5�F{���P���<�u�	��M�R�r�c���0�ϝ�����-b��Z)�49�c�B�R.M�.�.�~�I��`�#����
�K�d0�}�w%��d��;u?	kON��*�\R8u4�����a �����5�(ɋQlM�����_`�d�\̽��p�P�rw�"��a�ؤ�X�m�>S��d��V7
ɍ��dpO���,3����E�_A7�|�m���K�U�%欸��"�"]D8�'dW�w�B�6��4�4�v}~>�Y���>܂%�T=~�ϫ�7�����<�e��nk4��<<(�U�4����<�)���3��
=ۅ���],/�W:3�޻��&}n��%1�PY�I����)�-[��6��F÷��a0��?��_"�0=w\IF�K�@V�N�V� ��>��::�R� D�1�H������ݔ��1�ǣ���OG�W�:Hxc�"v%�=��jW�nQ�7A���;���Z9L)8y�W^s%˼�����W٧�ݽԚ'�g����'�K���d-��i]�+bzmk��j�V��3Lɗ�TϺ�Ͻ�/3x�<[%+���r���' ���uo�Km���0�Lb�Q����=�?z�Y�x�<NW�+�|��&����Y��K�L`�0y������%�{�����m�;�p�?0C$��kf�
`xQ?�"�D�L�z�����2�v�������4�N�~Iآ��3����|�S΋4HM�&G����ԻHf�DKw�"�Q��wỌB�-�Ѱ� Q�;���n�<�rnԑʠ�Z��d����"ƕS�ZQ��A?��/�Ś��^����� fv��E�-����
�Y�Y\A!*ߔc2�fh��\~��SV ����Ƚ��VΒd>���|�O/�^����M�"���*읹��1Q��P�ڱ!O�dYs�p.akj�� ��@�v���V`h�)>*�P�4v*���;U.2֯1�0��Qgu'��͢������@n�
�'�B��Hs��L��<n�Z㥪�g�2xeO�#)�%ފ-����:���S�+��2!�K�$�.�0�� ��`��+ �C���W4>g*#������O�:�$5����������j%��/�mG���䀮H�$�P�Gz���\*uP�uF_fn��l���g[e�߸�8��f��ˍ_�7w������R?ޱv�2��)	ajpt�SV�r6
^����0ဎϥ앖(ڦv�m!���k���R��1c{	�s�
ncR,���p|*yF��X��⯑�D_�wc��'Z�z��hp	���Ȗ�
��Ֆ��WD���m�Lb�̚���?�0هǛ��n�	�sf�j��p���E&P[dgLIC��C\BI�iA'&;�tl������O���!�o���5��|Z�ͫ%e�����>\nn�l�4�.?BЏ���k�6�]�i�����;��<hǄ�$j�?v�R(���%�(�����>�Q*Y���}��;1�~�
��WL~���g3���芮]����J>���?K�I3Œ����E��}{���P��l������'_���P̠�x����TL2�O���^�
.zn"�];#_Ƣ`K����Q�c%o��W�������A�U�?PS��"�|�1t��|\�@���o���
�j6qH	4Q�U��.��u�����05��5���H�/� �,yeIiy�W�/V�{Ɨ �M~��:}=�C���5��M3�/�9��#�=���i���\	�Bq��D�}�FB�0h�;=\�=�E�UL˕�"�=8�Aa+���n�p�����	\��-�d��b���~���#�Q/1Q���3Fj��'7�V�*�q�KT$b���C���(Y�^zxP�L�^�N�|S�������NwE�A�5F�]?�K��`MC��.��d6fN�尷߾�����y3�(��,��~J��[K%�To|B(n�S��3�9�I��KC�r���m[�O�GSQ����@������"���#��n�k�j324P��!�DҜ8얯�P%����P��,�T�an�\�B9�/��6�e��f�Pl�����X}ؤ,�Kf�sb�g�_
g?vVu���^���oX�����N�N��������\0J�vX�3�����t�{p�x��bߧ�����eI3
��3�B�|8V��n�,�C�V���XK�	k����s�if�^�5P���O�{l
����O���,�����|���L�a��-�o:����N��!I�,��l�.����\�z>�����($ߓ)��v�l��W��E�?-x��t�YTwà�zϞ7������N~@���s{�c	@�cá��r�8�bU����ǌ�b�-�DK�"��:�)ץ��"���b��Z;O9��m���m���o�y#�R8�8��sj*���k���@�P��>fщq�(��y�:���.����~M��Nù���ͨ�]3�e�˛c��Gh�p����oH�rx.k܂x�ϱ��k+o�V�_�f����h������g�����~6��}SdŵV����ܚ�d��3�R�P#������U��:�����DT�F�Eu3Wg_A��L��K>B }R���A����r�-�����Ũ���ܒk�ζ�%>��-���J~�n���dlS��@���VVķ��Bpς���ħ�IW��[�G��3�<*����J�M��r5{�V:��dxӉ^�uu�6�P_��J��pN2�h�<�ǃ/H�O�f:ъ���x�:�[Lj�'�ǀer���V/������8�RF�wʪ���C�/�����sg�mms�{�{>�'�K�ٗ���)ncJtb��*��h+˺�����ҍWh�Ȃ&�|P�k�>�������V?�u99N-U�B�*M�L
΅���kC����P� �`�;�_�sZw��iS�v�.[.'��yjh���V���k��57���VY��]��{�D|��X�%����9����p�Ǫ� �)2W��v�%Mnzg������ߧ�Cg�7��A_�=�Jqf ���#/���;�������惎����̋�ѪyS)1�|W=T*('�S�0��Z}�f�E���C�{g�	�&��{&�@��&�����@ˋD�w���?��7�qro"Rxu����v�b��!:���fB����+\�H�'�f;��
����(��+z%�Z���g��+u9^ݦ�LK,��j)ƍ�Ý>A=<�s4�m�:K�@�j&��VD���s�`�2����n壼W@Cܚ��&9�}t�m����������s��Ob�![0��ɶ��M�e�U��5��ο�6��Y�-<�^�4����22NV���������>��$�O'ŰM���*b��1��q��{L��L���;����E��ॾ�+5��[C�Zn���S�?;T�\�գ0���9uV�t�m��c�7�O�3ٛg���?p�r#�q`��B����o�y�$�D�Ԯss9���A�J�#^��k�/i�du.h�Ѥ	�Ł�>����Ʉh�8�2̇J��~k��Kq������rŧ[O���)�ȲX%#\_�V^P�A�0�8�
�6Z�bK��5��>^�?(�����(r��+(D�+�DR{b+��
<?��ܸU%s�V�'@E7q�K�Q���;N�hì]����aT��f�o�t͌b�Oݫ�Չ�~d�)�o�s�����Bs2{�y0�d[5���T�{�h鰤s���I�K >`������is��-D�6�͑uAa�K*7����*����q0�gJ?��;7~���F͚gd�av�b̪Ŷ��$����cbw1זA����ˑ2�m,�֘����/�-oY;mdh�~��v)#Q�D�������%U�[��t�N/�>�H�4?a9ͩ1[ڤk�^!H�ӗ��ҕ*hjϯ���	�s�w~?;%�����I%g���F�����Ј, S��T��X�2�xZ�X�9�yD�a�em	�཮��Q�@���DD���Em���M��F��m1Rn��oi7v 9?$Z���j7���I^2�򙦐|�|[֨����&	��)�#����ҊU�>��~��];�t2��DCC�+T����Egn�=�vx��������=y]~�2���0��f`�X��g���Ej��h�8�jA���ZD��PJ������Z��ݏ�򍊲W@�T� &J��W����Q��FS�Qb��e?�Tx�Q"	��a�m�����T6O�t/4�>~��f*�kRF�.����(�	�ɩ�S��9��]ă�ҷ���~
�ˁ���҃*�������ϝ/��v�qXG_�����Ӧ��"Db;SkvN˨�Z���JR�f	&)�9�"l?�.+������8�P9jݼ.Y*���J����K�VQɯ�[�K�-�I��U����Sc�vl��&�RU�O�:N8�R|���#1��B�ҕ����S<���WO�B�Ȃ�_��|VZ�s4RqG$�R38�̬�:�ET�z����_�h!�D�E?�c��(8��,�b|ר.?Ce��2��L�%p-j�7��(��m��nh?gT|��;��h:�"�V��V�)�*{	��{@荑�^d�Ql �{�\���}s�W�Ww|�~({T����P�1��Y�ȩ�b�Wh���d�LU(+��+��y�Yc��&ɿ��K=��9�fh�U�/��br&�n_��Nx����j[<3��V�7�}d���s��nQN���v�-f�d^�y�����8�Rr72�lA��A��"��[A��ajO\�O�A�w5����(��@�rO�zm9ʝj�PbBޑ���&#���8�:8��G���&��Ҫ��@�W���%��jsu+}���l����o9P��KQ�0"(�t�c�$�v�0-���->��z5-z4��v�Bt���-�#��fr���Y�3��Ex�44�.����7�|"�=+�D���3"X�ڕ�@'R~��?.{�n[R�j�9�dm�+���Mg�q�����{_oD�����H������8�J�9�ht�h�&�tmB�u�GUh�����8^u�cY��,R7�LSVf�6��\��?�7�*�2���RG}/�<�-Vs��c�s�KA��-#���!���:%�	��"�+�S=j��ܬA�n�����wb3���(����-C�jB��Ӕ(��S��<��Sˉ��:���;�cE3Ģ>aM2<ۆ�B�	�Qs�+��q~�}O�%!��ή}C���x���hԹ��}��M`�.���wh�c��E�F2��9�
9J��H�vbS���S�p����w�"
��9��.^�BC�?�h��bpg�{v26 ���9I����mf ���f:e�ҟxdժNӄ��Z�@Z?3���<��g�C� Ir��bqW��S�e���j'ISLP���;I�(�����Я��K�!;���U`��"V��Xݟe�fC�����X׈;�����c+�+y�(���,�Gό(Ş�����Qp�0z�eF�ݭ��j{��5�ɟ5���r��a����$�L�њ�qHT��P��)�]k-�VԚw��x�����m�M���;r3{��Ӕ��)�EQ�4��׋#ͱ.л�DF�"j��
�/�WFY�7Q׻�TU�hn�ru$�Ps�0ꤨ	,Gg�Yt̓G�}N�Av���Z�KK�H�?��|�N.Z���h@�o���BY��ZR6�[o}�d܊���h�b�����J7�t���G:W�1��"���'\���2�+v�Q���<�.m��'���N/�ٖ�����l`��P�����(=����B���
P�� �nl#��yyL9���C�4�9\��W'C	Q��(�r�Qx������Eމ鿋�}�#�2Lz��0V:f��O?��g�g��#�Ώ�~Θ]���ͲK�ˡ���=PEa�%��'h��l����j��FI<�^�kt$i��s^
�n:�GM��S��e���-%�{�2ޔ�U�,�5�ũs�M�����Ox��3�a�m.�>���UdQ]?S�7>�O�fH-�s,��ۙ��{
����E����Oۍ.ʊ��bKk�_,���Je�Y��˳��F�ĮP��PrʬU�W��Mk�L\�\������pN�V�k��D�a���!#2���ĨKa�-�C3��(Ϻ�GG��̟���y�d(��9�2��F���O��M.�(��/�����΁� P��'Ut���f>۲���s�;-���МY5L��D�G~Wukz���/UX�
P"��P"�N��ya�f����������y^�g���-7]`�!��l�ݙ驵]�drA�����I8�/�K��_2��|wѾW�h��h{�\s��� ��HOB�چw��-ub��噅x�J�	-L��h_��"Xrܦ�&�"��M��K�ލ=�'C*GV@&��ڊϬ���-g�{"��i
�^tM~s]P^�͐��*�h�fUxG���6��H"ڶ��=�f����`�zj<�,m.��7����3ê�%=�[�i���V�T,���ж�}6������ ��h��0{��� ����BZ�r-HW��␭��؉�(�M��=� �}y�����hF(�"�s))Yά|r:-�cϛ��uGu�a�T{J_�.|�_r��(թ۳}M����b��f��SA��ҺM�<��L�����S��|~m�+�4�[i�8�)$F����(��eO������,��A�*�d&��yc�3ȅ�Vư���f�-#�	ps$�g���`�\%}�Z�?*�WE&CO��~�j�H���*d(�|B���(���l"�>�g�� U���qÛQ{a��̒���B�c7����[)RۙiY�o²ft2wI�+'H��Y���1��{�}�Q�cU+/w�&�]9a�b���#6S�4��{!(g��(}0�+F�al�@҇<C�K�R�'���E�)T���?��V�	�^|8�6� ϭ�B?�pb��}$��y�D��U�+ ��P;�����B��j�#���S���̵��?G�OK�s][V�a�$�Q
��aˏjO�kw�n+�ڢQ��2���̊Y�>���:��t=�"Yo\+��DH�$+	]��o���u/���s7�2>:�j}��5�7o�'f��M��9(?u��n�+�1E_���*����u���t)a��|��T�	�y�h�>���s��!�RZ\ic[E@{�G�� �}��;�^0l�uoN���.�w�o:���>��NVb�NV��<z?cq��y�AQ���I��c�����߆3����0_f�A��$��쁾��t�����b�0V5� �lˏ�\���dؖǻ�h���C�z7�.�ph]�­M�ه�i�Y��R������dE�Эdض������e+�f��4�O?�}����EC}"� �g!�Eg�[���j�����<��݃3,u"t�f��3���C�s�#fM�⭭)�+�\���BܢwiI\ܼ��S��ND߈]�">ů�zh��s��a����8P��ӝ.����|bm��n��>I����	T�Q���a�>�8�5<�5as��v�zL�t�3U��&B��yd�Id׎�dp����Z�?:��
04w����ǥ"�缍��;]s�p��_���38_[ƌ���I�Ŝ�
%]���:3tUD�.ɩ��I<"ۢ��h�d>�$�$�����(CUB@ŀ~ xk�v����S?y��W�� �>�*n�j���F�%@�a��5��d ��s6tQP���8%�� �"SHf2T�"���oK?`��~Ru,ވ;�d�K�����U�*�U �j��޼y����6�k��H�J���:��'��v�($r*�I��K�/n���Ϫ�����6�6���U%\µ�ˑ>�y���x�~��|?���n�M��P��_��I^����N�2&���+!��-;�~��Ƽ�q��m?`"Պ=��	�U�1i�<Y�ڈXy�Mv$� ~��L{�^�27���_�p���Iʖ��j�褁��LJ��wZ��S�<
�#=i�<ś��YA���K˥!�d.i{۾j��ǥ��z�G1��Է@HD�Ȥ�ݹBbG��Ip+�����F�;;�z���"�'%wړ�&�l��_�MO�)�0ս�Z�/ �l���=��{&�PSh>U|��8�b���@t��R�yğf�Y˅��_�̚T�*��Y�3-8������?���R|��g��K�?������zD�U!�{ɱ��e�7���U��%2]�l��29����S��E���~X[:w��b�,殸}�2� ��m�0��0�Й��=H\���v�G7����a�+*A���T�T�>3QǢq �q�'W��4Q8��9_;��-,�kk�f�ĉ�-�#�I^���% �
ä����,�o&g�zbÖ�9�3�T�/��h�J���O�x�i�#���;����h�[<0.�-+$�z����z�>���<�(�_{���QYwsw��}�9ZӺp���dd�'�xܙ�ES	�h���&[,�D9�����)#®�5T�ؾB�im��o�<�X�*~���/�n���7TZ1����	�Yh؋K�j�d�h�Ѭ���oWk�GZ3Lu�`�j�ɞ|�����~hR�<����e���������/��!'%˚�e.!������=�r
�6��>�����#,�kn��?��H{װ�����3����ή.��6yYi�;�Q��"��Pee��8�?U�R"�	XQ8��aZ�@Q ��ũ���@x�­�;Q��ټW@���HN���e!d��	�0l�d�PI���BCO�ҟ!�y~4��+�z�xi~l�������of�u�����.'��y����Q�Gi���.�a�,�8-KYV��_�-���n]�(�G��Vv�������2mfM��]h������$ɋ�Sh�$�;��ԻT���2��3)	��LD�%V�ؒ2�x�T�#����n�n��!�8e�ۮ�'a�XJ�ooLט�5~��4̯���[튟�`��~8�߇T����e^�?��߅��ۦX	�Q�R[���(v�ض��d��pf4 i%�0�;A�<��B�f͓i�NR����N�R�FV��ځ+�pnr�yx:ݼP�69d�i�MxR���(`	�k����4�0����kHfea��s�('}:e��e��T���{��$��X�ye����0ѷ%H����<]|�~�7���у����c�*(�:# <m�]JhnZ!Vo�U�=�/����vE���+[n��lzrF�9�(�mCN���O�M�:�^��yhDq����E=H{y������o��o�Bɵi.�ʟ���䷚�o� �g�x�Ꮾ)�0?��+/��X�c�qwl�bI�%�O�l�q=�>�x����*��kUI����qJN�2>�~P<�{[u+�1'��R:]�50���/4��y&�㰿�J�.T�?�-
 �B��� M���}��ИR0�����ry2H��;�Q�} �3N�Dbf�s{���ek �����+	?v�q͇H�����VS|������+�݋��ZZ�� �G�G�g�OV�i��>N5�eE���wt�I����w%Ҍ������|���^���7z=*�����h�ۅ�(<��ޔJ�6~���>}l�}	<,�n<f�TG���LT���8�3���;��� ҇�g�/W�m�V�{̊��=�$ђJ���4�7��b��ڷV����۵߽�D����ݺ}�ap��"[}ꋃh:���"�e=Wύ��|�='֘ۮ왐�A\�}��@����A�JӮ�f��v�2����eoWp���tɝ�~1Ȥ9�ٖ�.��c05��zZ=h���d�:B�:�n�M�9^���E#J�>���UN��y��ז �x��
�t(KTT���Y�(�۪$����{��
!�Jv�%C�0;!Tם���T�(�zeՐ�C	G�����Moi��X	�͖���5�sc��n/Ϲ,G�W@p��5d������s�I�zA-�}zRo�����MPx:�������3gV�?����>k9;��3K.�N�Ϳ�u����4eS�atb�G��
�?\�ض��Ǯ�I;�?+T(�Z�YU��y�����A��]�:�y�Z�i��3�f ׽�QV;S�ͭ�½�iLKK��3�(R|Y��3ߘ���"�7�{�5�t���w��D��H��Y�cf�I��oQ�&��q����Q��E��O�sU��{>��S����j�J���;3H�u'��>� ��d�j��Ԅ`w�O�"�R�n���\�����0�|��&����m��"'�7���:������O8
���i^��-�#����C�"��p��'A�Ѧ����vM2:!_+/}�g��U���Z���}P�g:��&kc���=%�X�I��-������:�sJ�������Ř1�?G��(�.{�#@��W����X߭�bN+i|����Yh��)-�LAO���'�/v�2��n9q^��lд��<�}.5eӒ��\	�C��1��V�5�2��W��ҿ>���h�g�8)恉� ��SJ
�D kF{�+`���N��='W&CP���h;p�B�\��M/��WM�_�$+�5AEx�b�t;��1w�_QpQ��A��.�Db��;�N�niA����n�F��.Jb�!���Y���<_ϧ���g���������$-ch�<x�7�1�K\(�g��_mr,�o59<]�k`d=��l�������n����8~�yzTXt��s8ղ)'�-.�����ë5u%��Ib��+.�Z;��b�;�G���ފt�������C���F��W������H�$�A�-n���q(������3{2u��$	�

i݋$�A�w�F�?d�'G�<=��m���;-�M�,@�AUt[;�'ҭ����6i���{#Y���9��e���ц�ρ�.3ҏ��X��q��b���+����	q^D���/���z��|��{��dJ��v��֖�,Vė"A��lK���Ja:JO%V���8��ei5+�>�8:��d�#�E4�G�����?!lʄ��/3�_�7�^�����FQ �*?���&X��'��"w�9�o��"�4O�m��S-(�ۋ���9eWm�C�,�����cUA'��kL֏)U
�� m�;�jڂ+S3g9c�v�h��"��~J���1/��^�l�n�ss:~��K�ӑZ*�WHw�� �X	�ˍ/��f��T���EƦlI�2�)y��h��C��z?t��|iY�%Qa�} ���5�bW1��'#ܐ�<�@�s6�5�۰���c��"^��^��8sj��Т��QOV�m&_��qכT,if�(�t|���Ř��zzL,��5�$ϕ;k�<��v� ,��9d=���/ /�dp#�F�[XI��;ĕ��Mxαq���@Q��Ƨ�y��|p�;k.�g��0�9>�����!Lx���I�F/Y���^�櫆%m��M��p1�3O	[H*�����pr�Y
~���g�$���Q"v-�G��Q���cϞVz��~�\:f��4]{����Y?q���Z�SN���K������h��cphRv���/���S��/3�ⶍ��T������bk�r�1�G��6��2!y��o�o�zۆvM���W��\���N������$b����vySD�nuO?޷�܄�4|L��Cr�|M��?���Ѳ'Ό'O��FH֜t���;�?-ˣ٢a�Ƞw<���Bso�j.@��z���O-S7$;��X�)*g�r#�$�� f���� 5�&ׁ�^�0@��*(�F~���/�q<�*�^ج�Bh�#2(�흆<Zw���֙�7B�m���|]��d�8(�P"����m�o���ʕ���_��j�ͭ��z3[�J��`VS!yC��R5�����Ynn���|x��MR�3{J�?%�����T}�~wy�D�����W�����k?�'�|c���S�%�A�u�<Ϥ�l9[���;�P���Y�;�]ƈ@u�z ��y�L6�I9���}y҄N��bP��isS][�����w_�/��()�]Z&�j{�s	��[@��@_ ��vvV���X#
�������'�n�v$��5$�r�f.�`�����V�ɇ׊��E�*χ�+ds���:�0�uEs<�2ޣ��uo6|P�<Pq+��QKK`�"!1'�!o~�-���P�K��GF�ᐪ��l�K�X�'��d�J����(��1��?�Ԃ������ �lA5��$�
%O�v�
��T).2�T懼2�;!~�|T�5D]ۭ���פ!_�����i�]O�	%Ϯ�X-A~��h�ߪf����������>����~�tAIF!wRW�!X��c���n�cQ���/(�A�܎`3v|RE٪ߴ��G�ϛq����tu�����)ch�:�O3]��{.WWp�jK���^i��Y�k�Lh�e��yHz�W\Z�+�1!��Q���V�wk�yKUKy���w��:T*�jt�&Ne!�V��}ˋ���*$��]����N�#v�Ei��I9J�	P����w�/��M���
x5ճ<��Eahg���S�?;γ�Co�;�ą�?3���c(b�*ǳyX/��R�O��|�:8�Cg��h2���  ��^���i�Y$�9�+ut2�NF���2/ y�ǿNn���&���9��
;R��8�06�+�މ�W��3NŇGN��AW��/EӾM���h���?�%��Nߌ�徤I2֮6k�O$�V�*��>2�>������[�&�L��`?x�v����9N������7��"I�~�/���{� �/��T�ẃ�+"_L��碖QA�j�g;QĹ��#v\wA��{��^ټ��.�#I�^�Vk���Yh#�[������Q �������pc�>H~㠛��J#���z�Pz�'"�6�Y���I�w.SB�;3|�d�gm��v������vq\&�����1��h��W�(��99K��;��&�l�����-l{R�` �Z�o$�v���l����	R��xU���i��������sY!o&` ���tZ�8�]v<��[�4��,�ȃ�͆s��F1�������������{�e�;´b�T;U^ 1��v�A3��gT�lo�ܨD7��&�9����E�]���4X渰}|cU���/ �,X����!��`��O��;���� ���&��k�����h�d�|ìf�y�Ii˾�^X�;��.<1�
�j��\ .�t��c3����D-�F,ݔ����j��)�����BY��׆�%9]z��x��/�JE	������2 �T�Y�b����Ԡ����qe0vϼ���@�j�;�l�������'}yw4���J�`�+B�&��W��<��th�$�xX.|R2L��u�/Hʭ�SK_>
�֪8�z��ڪ���j�z��6���k}����Ln�t�X e� ��^z��X��@�ƒj�A�g�i�[K}~rTw��+��^8LDg@�8���JE��Ga��Q�m.��J��E�\�CCU��ZΒ�2'��?���E�\��	���*�GxW��o�W�4b�s٨uS_ ��"Z1���-4��qN�l��\�{�2^�\؆Љ�c`]�f`fr�~�Ĺ�F����>8�^��^&�Z�
�a��uޕs��d��j_�aF�/ Z<��p"r[���ٟ�9���f�/�-N[�$�>l�J 
�]�ӭ�Cy'<FۼӁ��s[���-���J�
��h+睴	3�CZ\��Vզ^�4�?2�5LE���b�-v�>�-��K�?C�SM,�S˰�lX�	i�Ͳ#��nGSK��+ ��wK񉱖l+Rr9T+��4�������K��=��*�\��eYE��SĿ���!��s� �5��SS� *��Q9<޷���)�DV�<��R�-�/� ��5�ޛ�߰�$����m#���܆yE���I��	榎�릟MwND��do\=?�S�O��GCg��\a�b��X)���!�^�ϋ4S:N*����g$��2���A.�{�x@���f�Տ��
d�l�ltaO���x��e�+��	X�S����>�ǰ�tμA��F�i�[�e��-�?��^��I�u+Z'97uR�ßk)�y�?  xΦ"E��i��k�Rr���[�)����0�g_�ِ��Y�ľ�Ί��I窚�Rrqm���2�4,bR~b*=�˩[j�q�A���ݱ2U��	�}R�P]Q�k���M��K`��N,~T39��	�^��D&j����\�2Ї�����M��4�I��SB���L��u�'��:���^���عe(d��II^�_�׃Y�^ ��u�a�3�V��G���R~b���kD��B�y¥v4�U1	YSr3�i��T7�`���&�;Cv�����$�1�c�5a��yy�F��S�����ІUk4A��M��j-b�������+p���65~j	/�C�~[G�������ns��eR�����=�tps'޻U��խ]�ͥ�uo�p��Q����{��~�+�2��-�3�]"�\�%i���\.���!W*@8c���1� [p,J;�c֧oi���NH,�Q�h���DK�	��/1��q? ̷�	n���J�}�{�a	%��Bb����:����=����ăȚLf���.Nm�ݎ��sD쟾��('�8�U@��¾�^9�4]�{m�C��j!���Â4zLN��̬�k������'�@�!o����Mcmb(���Y��R̥�{���[��'~��쭎�_�B����3�/P�禶u�J�SR==�u�ْ��HY���[ӹ��W
�,�4K��	�i���fo��A�r+�'��Nލ,��
uI����3�+y�z����|�rg�/�6L	��jX�%�y,]y�LQK��H�H����M|g��s�V��f��Q|��f�%��]N]^W�I��G��|�OT�{/ lo�wjf�����BT<qΎ2��М�ɞ��^N���})�O	i�E��U��+�#�w�M�ՠ����`��r�-�R�[��)�Ry/m_^w�4�c�$���xՖ���*���7I_9&�n6Ҷ$9.��� Ql�jezvD�����@`Wt��$� l�M���>�몘h�9�3����^tSl��^]~��&�2� ����pS7��"F)��e�W�����I]��m��[���'��Ƞ���K}u����1m�|�d#(��?JK4�
�z;�߾�����"AK��/�W��<Z ��\]�������ԍc�8r�B�NIIei���Iy(�`���x���|�y���C�`��PmJ*F|ѯ�A�͒/�ox�=eOSۛ��R�6� ���5��t�j�BJ-N��sd���[���j�А�%"��2NM���۝$�.L�2N����-�7�t�~�ӄ9\����h����J�$�v�I3�̏Ѿ=Os}X<�o�%8�"�J��Q�o��ʒy�ª�Ѯg�+A�6�`���T)������-O��V��S�L�P����-D �0��]ʺց��Y���(b�=�}0??����G�����9=���rU]k�m����C��e(�7J�L�8�'���C|L��v��-;��z�>E���}ۢ�.R�.wo?#�֘�$qP���^Eʭ��Ԍ���-�%9^���$���~:u���%�ޥ<h�m��{�>:U!:��u��by���=��<��uy�o�^�/�'�t��mH�����^�z�F������[�ʽ�p��U�<�P����R1�ݮS��c�f�+���;^&q���%T����4����w��e�3ٱv���uډ�fʫ���u�g���?�}G�a���ֱ�1��'y0�+��!}��Bnd/�ym�Њx2D^(Ğt��,����0���E� M�_�
�ZNiV�rï�ZG��=��_f�FLͶx��]��>��<�$?/��)#�}�'�
�k�||�^��&;xOo���"���o�XJ=��ɭ�"�)-�g��,�P��yvA������R�������W�sMys��Q��E� N+����߆�q�����~K���Ù��{	���(w�Q+ukHZn/?�s�0�):���t��iV�X�Nгt=��ʱl�S�("/�"m{��\�N,$��;��QOM̕�ZX^�\4�x~��6J[_���潙e��M�\�l�	��.[���i�q�M�t��M�x�S[v��(W�J�'J�^��y��>����G�"%׹Ufe�v��x*��"h�l��:��}���5���vM`�x��:�L���_K
=��?�&��c��&�j`�7z�sK�v��~r􌦵�F8���)�el�)������%�&���]3���zl�4�ʪ��2��C�to^����%
ض���ϣ���~sL�{�#x�?��@�]�8/`�./U>}�'F�6Mm��B���G�~'�~���K�
wY���bX̳yP�y,�0�]�y-�[ױ5GF=�����U��A�� A�P>2o���ؼ�����?��仰��j�l�jf��A{C��T-���p<k�cT���ў��g4A2��[?�V]���%�(���p	6;lg
	��@���Y04�Q0"��'1x��E8�Ф�p��墤��ybᆫ��y��b�~�]���'��n����M�h�qU684
����̃�R�*$�
X�)��NY�r#S�ld�<��{Y&�T�����ȷ^s84��M���;�������w@�=Lj�v�-�MmN�v�Z���������8�Y����R!�a%�;7#_���'.H*~���Yp��L��^��M��2�R�c�����睈��	��Wr�<��G4UfH���7v��+J��P��6Pt�/�6�D�n���dIY�2j�2d?�����tu��>���1K��a]#�ڬXՔ$�B��
�,ޜg�q�����.�V$P�𼓡euU��4�-`>�p�l
��A�7	2f[z_����dʩ�Ey��^}s��q�<*ӂs7��f�!������{����=�vB�~_��K~A��g�bc2�G�_�kY�?1=S����Mp߿�R�])����N�=+��x�����~��ۧ��99v������A�Ż\Q�z]#e6��(�8�|L�_ߧ��0k%��?t.�y��s��*��9<�(6���
ֵfN�D�G&�i�`p�2r3��p,n��WB���Ԛ�&���O:"���\K�̼�1�Xc�Љ�OLp��@E���&�q�Uu�}���x��l����-��9E��A33y̐��FpW��/U8��{�VZ�F]I���pʹ�
��	��'TC�;\����<� 0F�κ�_ �_{wӄgx�a3�(�C�As�r���z�Md7��"adn�%�"�`��{����Ն�%�3��ռ��Dkzx������h*����y8����i�s;�1�6�_�<{�vF��^��3ws��4 ��9�N�dݳG}cYl��zgl�|ט0on�=��=�6|"�F�J�U^i_aa%�\U����&��	�D����fi�{������hCUؿ�����tlA�̻�`��r<�f�N�IE~:?I�Cgu*��L�H1#�G)[vz�:���H��<L�i���PF���(c����qT��L�>�i�N�IZ��ظ���a���D�̏�}Ļ��K��� UTR����&��<M�>D���:9Nu�F���!��+��B/���:������yu�R�0���K���ܠf+����$8�+�}Cn�P
��*F�B��^:� ���_ 5g����?6�vp��%�/[�{��ZqK�2�G���(���;�sEJ���7ŉG�;�3^őr���&�N>��+#�ǟ���Y��yo�"���l�kC.~�S�ߐ�����v>����jSu.��K����D,�6fWb{��i���	�T�=�����OԎ��S��
��fVD���������,,��`���U�P�����Bl�����;�S��x��|�Ąg�`�����2S v����[9�b�Y�����-�P�_C�y�e֘�S)G-��+P$l���g��\�esxktU������w��w>�ۏ�DɭR�,H����|��D%=t�Ha;@
�r�떮dS[��zG<�����N�A2��igyK��&�p-y�����p�`��v1e��Ր<�i{�]�������~［�J����[|_ 6���(���0���8���E��u������Q>�����������9����`�Ψ�p�ⳁl �ߡ���FA����"zM���4ӵ�v7�ym��X����y�Ss���};RT��ƾ�>{3��â�s�Y��b�j�_�o�o�LY�d�P���}IҮ�*�t/ v��5ٓ
OJ]F8<7�aHm��Yn�)��Ť��>��-�C�+�.�c�	�Tpꙉ��p�R4����l$x�!]��A::�����]SB6	�ǡ�����{R֫�ߌ���Ψ����}��I,�.=2�T�b|�e�i1S[$&3r倆��_��SծZs���+��u9B���_m�~<���v�/��Y����D'����G��o�!Jx���o�&�Vڗ:=�]0�7����|c	d�>�a�)�¬��H�Z2;ZL�:��$��.$`����s�Od��ޯP�G6�K�1n4���.�4;Y\��n�!V��'͆ ^�5�lC�`r��9�u)=�*JJj<� 
���!ׅE��ךs%,��χ:��?���r�ؘ�h���W�A�!���e��Kpk�idb��Q#&�����g��$[O���rGc�~f��S�։���^��i���`��!d�@ø'0��vnd�(�&np �X�g���¦�B���K���2$�����q�난D����6�<�&)β�gze�K9ɤ����eA��5;��[���E���`�Ȩ�/_�q��Xf�~:q��8~N��t&���V�(�VV��1LU�"s\��d��ǥ��&=�{s����_��̣��5w�T���$�.�>4��R�&Z/ușt�@����}�<6�{j������-hO���Ñ~T�(��ؕ�նc:d�jq���^�
��&�r�ף.� �E�Ao���:	�h���8����;���.,]5����"����z�ֳ�9�yU*bʉCy�	��X�[�^.�ls��j��}34i�_��K����D2m���ϊ�� �P��3�Í����sR1��a���
,ienmW10�/�汈e�;\��z'DW.��4�UasF�Ԝf�'볱(�o��`JoZ@��v(�x��술�@����O)�栧����Z�&�7v�}�X�N���_?�
(��z�F�g��+="C�q�/2���~�_߆�݌��C%w�G������j{묾67���JL��bh^�?q�����  ��C3Y�oPa��zt~�
-$�~;:� sd�$u��^�GUfǁ8+_��?J�wy_�\� ���q�R� Z��(=�����y�g'��0���a���{]O���4dT���X�I�f��%���e��Oɉ�y\�Y����(С���<
����?j��R����("
�wC8��I�k6���0��P��3�"���u���{����	�K��V/���*��V�m��#V���F�T2}�yTq#��j@JY͵9��A�?&VTp�L}��q[<6��K��{ю0���v��h,�jp[�+_ݢrM1�K"��!ɾc��Hi�/�ݏoe�O���v�p�=qr\wШFM��˥�q�r?��G����D�m�bV��a#�g\<y<����#S�������h�1oP�����"�Ҵ5h��<�&riih�R+X% C� �:�[Rv��S��j� q7���|j��\�j�|��`�T���}~$��w��מjcs#�����e��Q��"�p$з#���c�D��E�G�-aUS�v����Ym�O�j��9!"�V!�@�!	��]�OJ�~5��������ֈ�%f�����!,�%�2L�
t%x��j�:��&!]��G�vvj�ͣ���әw(�o.|��`���g��	O�y�eȮ)��&���;V������::)�on���d�gn�s�x��[��@^�d���Kq��$%�O��p���Xa�����3�d-�eB~ǣ�a��[[��E���s��ZB����`8���$}n�ԓ�����ҵ��!���T�^���!�ni�n�*��\�V�q�����z�2QU��N*Ԉ��z��1]�CFBq^���Y�{���g��?�9ޯ��u�UuN1�d��`�J=�Q���q�[��6����8"�@#*xRJ�����}{,���uE�خ�M&.���aĸ֤TB�O�1n*/O��-E�����\��z ��	si�U�|�*��Ш����_���'�� �UGg�����U��\G�B|�r�b��NF�Q�g�2̣�;�/魅Aw㾨���y�A7J�W@�#ӈ�H������ɵ⥈7�t�$c��̿	��P��f��Չ�8�l�%R6룇/纭�c����6��Z�{HU�F1��<��z��n :��y��F��[z6����y�<ٍ�n>r2Fn�1Kt��iQ���<�l���@��H�Y�Y^�
�Fq"������/eC�7
��*��ۘ�N���֋G�ASܷڤ5���g�|˂�7�N�WLr�~�|u�¨���n4�C����4֛䅍�Z���C�GQ�Gz*��}���y�`/�X�Vi^��f�H��s��@�(=��g�"ݣ��+*��/ l��jc��ī��}��6Wg���r�1�5��l_3T^hiV�";Lx�8>ͅ��B�u_s�����f�v匹��QS��p��=׫�+߮�;+���	����#�u	':��Z�kd���(d� 	h�w�i{�t�Hș��;�:��UIL\���}�'��\e�/ �oRH�m�7%�N����`4��ĴJ�Ļ�AȂ����O�<��M�c��|�W.7/ �3�xm5
l9�:�maI���$�sc}��䩩s���1������v{f�ߋ�o}ۘ��h�j����c�SΧ���x��.~>��!x=|}vzc܎�=_O�$s��x(bˣFJ����!�e�������̿m�@7�͍�h©B>�.��8�:Q����:Wjx����	��w}.u*����:H)&H�@o�t�\T&ͳ�4+G����۠��� Tgꔄ���슴P���1j�+����|�&�e�^ C��%Q% ���ɺA>�K��w����4��������و���rM̱n�^���x.��ͻT>c`�;ؿ���U,�6�b�I�K#�g�ʎ�)�OC}�����\����r]��М�Xu:yc*�fh�-l���/"2��	�e��ɣbr�`������<��	���i�����7�@u`�\�B�����B�k*��c+�K��^ �	N|���N�����t�;`r�kM��i	QKE,g?��OFc��d�gJ^<��r��k=�ZD��{d_�h�-�k�'0�'L~���N{����i!|��� >�.�` z�x(���p�4,WZ(_f�JF�K�a��4�&A���Jl���F�����B��De.�`��ލ���;����-*B_�G2�'<8��%B��Y�f($A�`�M����ӧ�L>���%F/��';�~!;u9_���;zz�D���AT{��Nb���o�U���y]�h���I�ی����Xc��cӡ�W�V��W��(([��\>ghݼ�
)�,�W���� �Ѥ�j�F�Ƙ������R�Α-�,��&a�pM�9���ɏ�
{�^�y���ȵ�������3	|ם-N|�7�[��|ح���l���(.6]���Q�"����C�J��Xgn��K��+K��S
]��n?6�LȫU=B���#���ӕ����{�	��C�����Ȟ�<��a�s'�n_�X�r(��[t���� I�h"aAy��%�F�'z%�&�cdQ-�:��f�`�(~r1G�3A��|T����y 1)k�����1�$�����:�q��ϗ�D����K��[J����? 
-�)�!�0_/W�1)σ�[�Z�~�N�X�0OǟT`M�����]!o����t�H�w4�6G�%.�Z����&(��`^�N�f������td���l�)��A��̊|�����G���oU����(��<�:y��ZF��@S��XL�,!T�*�� +���49|?Sz�M�n��9{��^E���9�n�ei3��&N��Z�d�6E"��,Ȧ�<���7H�W@(G�y�@��Ӟ����F�@����� ũ��
���TX��6>+�0��'��Y�s�tB[��D��x�$�^���+��#Q�;n��RĘF�W���X|��X���ˊ�|$���1d�<�&y�R� �����샳�슓��-��x�>X�d��n�#�Z<�V�8~kؑ3��-*�\���\U���)�(����3e�ũ��3v����������jS��.����w&������p�D�$q�
;��4sM�`��L�:��ӻ�_!<�>�H!=�P=�W����W�C�)�6:Lx�rgB�_��и�)�W2�M����b���~��$7p϶1iH�c�V���:wٜ!����2�hU'��c�-������]��}�P�81��N]��u�3u�_��~�<#��D#�|�6��F�ٱ��iw�z� g5�q�w�g�rH\/ ���N�@M�*�<�f�!���u��	���2U6�`�����b�����U�k,�2wy���m��C�{u?63?���<����Cd}ҩ:o�f�����C���*��f	CǙ�Vq��D�b_���KYN"�.!���yK����@�x#�m���rhG����� uc�;l�D���-7�5I\��B[��r1{���J�0o4�1u�ƀ��C F�z�ɏ��p��>�g����l�[c��M�Ɇ�܈�}�R����Q��ro�`��jw���ƾ��.v,-�� ����1�SkV�^��@<a+񍷺��Bea����R��$�����mG[oеF6�nQۨ����k�D"�� /X(iK��&e!ן����������JY�K��'t��jP�V&�*�D��~u9s��:uN[3J/��O%� H��Р1.�oD�%_ZA4�!U��849�^�%>IWãMS���G�vv-�ڒ�?ΎU�
e���ʀe�M9F�;+���>b��&�!8���D&k}�5���̓�@u���X�˽�T+�g���M��?�P��'a� @c��i����a����{a�C�<IQ%񧅆���?�SN-L�gs[�O0�R��0xj���&�g���EjM/�Uvi�'����QakP���\�E�G�7F��J�ab��x7FX����Ξ{��a}��;y���"D]�hHd���h�K˽g�sF��{K�KϹ!��_�"Ĵ�R���r�L��9x�uZ�Uo[����s���Hg�ʭ��I�D�!
&�!����'jz�h�y���4׈��e�i2w"�Ej�K��Ʒ������	�p�YV��\ݘ"������yiGc5>@P���IDY�_��:C�>�g��׾!|�����5��UI�{��Dt��P�MaTٽF]vo����� ��{��E�Ձ���E,O󮓧�~�Cy�^�ܟRyc���dA����E��B���+ҧ H�)};���mDXNO�V�u�v�uG�qZJ�g�W���d���ȉ+d�?�l�yaP�_#6�P-ŋ�g<pJ���!�,�]���e(1a��@W/fJr��bA_��*q����Ȳ�_�����?b�xc1�j���ƬV���ڒ1�+�Y/
��2�5�ښn}�)u����+���>���[�C���Hn�t.S���#r ����_���Zc�iyE��!�\|,(��S`D-�MΜ�����L{�<}�;o��"����_�ch�V��j�V���vJW�Q��K[l�9�fzrj���ߜ%f�%Pl�h%�޸VHvqC���sm���׽�gxֆ�odZ��a�}�ٔ�U���,/M
�iU��ԋ��/+*�u%Mr���DY���
��-&�D�CB�VO	�0�G)�.�;V~&5y�܏8i���R����
�{���IB�*k��2B���h!փ/ 5�֊�qM�5X`Z�
r�#�3]D��'��Ӣ3�t "���=I�:3Vh\,c5�dV�`�^0� �g�x�F�is݋�����t���;%66d���������W�M�C�e� ފM#8�b۳c׬���ץ��Pఛ�)�{����.��$b��WlwTS�LN~>e��Q#�<�>�-����_�L���l/� �z\^�;�}�b��99�9�;~A��b*���ǑhP�f�뒷��e�����4������M{_ˉ#�O^�����J����v/pC|����ɂ����L���&?���L��O6�����z_�_
���?��^��kk�h���I���wQ@�+o���s�����B�$��^Y�"���)z{���[?�#?"��B��k�xУ��^�����蹋��п]!L����ao�sU���3�̙�_I4&A!d���
��4FxI�b�+���(��q�l����D*x\6�5����� ��1UU���t��3ߏ1�z�֧i%_K���F!�Zn��*t1+b"S�ono.��������K]++��h�� ^�\N90�k���G*/�8)�B�bk�M��v�͏��c����H����&��f:͚��,"������ņ���"$&��d���I
�"k��H�i��e��8Y[��h�R{��T�1�'������2����y�E���չ�g%1��4��@9G5S�/G�ڼ#ܫJo�ه�1~qXwoC��%/F5�� �aa|Z���Ycb�^���,���U8���	�J�e��=)!��"~*D�̳�/ 4A2�G���U�Ν�!]Y��-�x&#�Ԑ�RV�w��%Siw�4j���yD�^o\�~*Y���^=�����7u �����>P�#���U܆�R�-͝�	�U}���wb��F��A} �\�F���C-��ͧ����|u�.4}�ɮ�����[
q\����ܯ�<[-��m��
����ZXb�4�g8��������w��8�QuֿQ���&��˯��zB��k��W$mmw��*����7��74�8N��1vPz�
��#��a	�x���W���U;��h�����%�/�zݧ�s��i6��1-1M啉�:��o�?���o�����3 ؾI�=ӧf-of����;����k#Ô�L������Qȃ��䅍��z���jީ��u���>�x
�eo�F:I���7/�?����k���j*VQaa�H�|H��7��F��͞�iތz�Iis
�����k�"���*�j����8t�z�V1N��K�=�c\�v9u�;�&3��m�g$�%�\�@��v ���^��!0�W��I/V����N�WXn���ϗ���M��Ym?��*���}t}��|��h�{N��N�����ҝ+��r�h��+�b����Ϙ_�(�d��a �jH��Q�ǽ�K�1��io���oں3��T�*E!�i�@��z�\���2B�I�fubm��C�<?#��(�d��T��T)w������}��$3��t_��oԈ�]��_��˭Jr�!#v2Q�N�K�T��U�D^_���(=��3��\T�}S��0�,��{r-0M�.ˑ����w��Vڌ�dP�?P1-�c8�)Ә8�,>�KW�mZZ����Jy�IQl>U|�3. �J��(�FYx�a��{�$��c s ϻ�����o
���3��̹܎q}���?�:H��_������m a��!���RTdV
�ª�fnmC��j�T�='G�h�V#�إ����Le]<H�iّPt��'"R�P�צ��Zb;�&�X���C^��DEȥG�,v�y���o�]-��2����3������;{D���$�&�v[ȭ'���܊j�ep�v�b�ғZ�ro*����$Ph����_F61Vβ�Y@z@q�:,�E:�~v:��FAp��V�_C9��uS3��iI��i�MFW��1�,�����j3|P�C_�&3;z�;����F6;@k������k�)?����lM$��?#+'���5�M�ח{����o�+��%����*�)	`K�Z����ShN���g�9L۫���Ak���3,�͹=An�i�����o���鷜�ngj�'��oh�A�E9���}�]!:��i%ve�u�Y�3��^7	�-�z�� ���]�hn�?��b&4�r������x|�j��VSf?K���O����Ys��k��$j���Zz��ߟ:����G�n��O)u=�u| y�k�pp� ��~P����b�R`��� ����6�Re��.P���%��>�[N"֥�4����*{V$F�m�x�o�Lo�1��8�1+�bs����3��"a�M���1G&�D�U�ň7P��~'#�Y�3��Xn��wc8��D��o�������囧�~�Vc*�T�g>���v{��c��S�\���ˣUfu�4S�\�%&(S�DL���쓑+K��@�jා�ք�6GO���w����GiT�B_ _���,^ O�E�)����p�ߓ(A��(u�[��c��q+��w@ ���7>nZ�j�+f�m�����-I��o���(f���K��J-Ne���̝U[M�n�`���`�	����n�!����3��%������v޽�����>����zz�z��/]��#��ݾj�ö���(ݻ)�jA܏�:B���[z��F�I��t~�͔8�-/x��t����i}V&n�d��Ϗ�󝨺Vl���P�-��IΑ��ߞJ�yNl2`�0��#F�E �4+o S�W���\r>�����kZ��(&���ׯZ^���l�tQ��i����4�靰.-I_45I�	
�|ͬú�8]h�C�Yؠ��ũ�!���]�k��
�Z}w<',+W~��g.������3��-O�O��'��z���]��v�u�����y�����KՂ~5������2m����.#q�:���\;�c,e�@����z�qO��߿�t���e�d�{ݯ���r�pr��gdvqY���P{��߂�jv�=����㇌���zܗr���h �P#/�%r���=�=�v�5h���q�)\
x�Vۙ���$�w���UC�DD���Se����֞���RC�!���n��zI���wu�8�`������CR��\;}�$RW�6����{�Hz�i`�O��ܸ���R_-��j�=^�Lrh��F��T�V�h2�^�p���`�H��K7g!�
�z���m�1��f�]�T��2���*,��G� �tP�R"���)nh��;M1���yc� ON+����i<��֟��C�N��R�$:�,���*x��F+[�f%�n!m?8j*�1���<�/��G�J~][-ha���#����/����Do��BG���x��@���`<�@
���/�8۷����_FU��CL[$_��L���|�'�Jb��xB�d%�uw����)��Fx�D�q��J�m��
�sE�as���¶{�7@�E�cR���m�N;cC�}e��K��*c�bjc���&�XO�A��..Jsghľ�CXw�2N�@W�S����9�Y��,-�'&����^\��q m-\;�ӳ��~A*Κ���8r���� xG��>�z[�xy�;T}IK�����q�:B�S��ҳ��(��A��#.V|�%/^��4wEB���6ؓ��,c�˸!	���/JL���X���Oյ�MQ���GF��aa�G�۷kТ��W8 qڻꙓIa��ᨩ�p�=	=Ei�[��c�Ob/-5"F���8�zyi(,`dr���s�iNͥrrk�����LΚ���F=����
{߅��p��l3�wҾۍb8��q�z7�/ϫ���O-�qP�A%��~:oxz�6#=v�pc�����(
�9����=��~z:6��b�X[]��|p�p���}0��L݄�	G��+(�����c���eg��7�ç]\�oL��+@o f��O:�x���hÿM��@w��0NݞQ��"7<�����1��H>[ /��%.�?��ᒫ0�V<��/���)����t?f`�q��2AT�ޭ�0�o]����af~Q!eC��A���YA	�q9ω�o����%�x�yU����$E��~,��*�����OD�]�*E����@��(�ڂ��f�t��g�E���15�+����cn"Q���A<����b���[K�4�F=�+��$t>�ȶ���������焩|��b�+)�u��o��Z���QHH ��g1��+�i�X�Gh�J�*�P�s������ަX��|{I;<�7��_�1����"F�R�xcXz?JTV$ۻ{��f⓳in%��܃2��2\����_�D��^���e�m��_�{cw���bM�9WRz�/�x�m�L�6J���틕ל�Y���O3���}b��]� Y3nv�s�.c�w�1�hjA�?oj}�ux��Ki����EZ�_���iKd��RO��/9�6:}������w�]���q%���!�<���Q�A��ǐ���|����KyJ���+�����>w��m�	��˳�dm
;S���!��gR�:��������1�T�p[S���e��Cs�4�
��R���v��M��#�J��?�<�Ͽ�1����<bO��C��p?_�Y��1ܞ�?�"�O��ۭ�JWƴ��+Y���[��$���!�Kr\ �����f��o ��-O��*I-�~Z!�X����~�X�u��{r��Aሺ���2fK�B!�3�U�<��^N�ENi�Wzz;z���v�"��W�t}���"[J�q�)���XD� �����Ӓ(�����D��ke�9�Q�����/��mQ��0������Q�,�xH���|6>u�h.��2�i�P�R�/����٬Y��-�l0��:w^�&�:ޜ<i��o���z�����ז8���gUc�=��1���١��o��ȍ��=��!�3�+���0�){��L�-��	m_8��5�*֟����=����9���������x2{B��7,����@L����1��O�/��P�S���r܊���$J���=�=yr���泌�=&���A���F�'�����n�&��׿�j$�1�`�fz��D0uZ����;Co�!J��> sI��_�mDl޿(lַ���Q� m�����w9֤�����q��?Ո}����ny�̑2�2��99��֌'IEx+f����xQ1z2�M��+F�M"p�|�n�[���&�s��u���p�웖�~ec6�҈U9։.�}Q��A����0r�E�jpKj����yKҴЖ���dD�|���?�$��m�c��8+3��4a7��Sg�`(��Ε�54O�����_ƈ���`�O�=s~6[�?������n���cvXH@iP�33��L�I�g��M��M
!�����C�V�����,�V�`�7Q/u9޿� �,"|�i��{$Ǽ6�=�k���ƍ*��DLF+���a�/��P��������︞sKV���hI���(.t���l��Qhd$Ζ�B���:Q���ὣ~��`n��{��P����R��`���w2\��0T�}S�&ҒR��`AV����m��/�m1ǫ���
v���ͺ�����8�~>ƒ�z�s ���q���P_�Z�"�����
�.��=%���x䋾���]7=#c8�U�]5�?]s���i��PC�ae���¿��G��X�c�����/�F�=��z�%Ѯ]M=�Ӗ��i�յ+�p��C����P^RJL�lH�%��V��O:!�]7��Z���.+pHO��fO�����o?��I��ӶQ|-'4g��bt�u)�a~bQ[%� ���E�g����+Q�gYιbqvW>���NV������YD���E�����Zh��D�	�'�k�T/�l|�X�L��{����|��`����_��J�{��h�׺]4n~�חq��0� \Q����;jV��pŇ�Ӗ=y�	�X��>GS>a���6ח��,X��AP���$m�l���<�#�S���#O�u��덃��K5Jz�Ҥ�O�	X&�$=��e'y�>���,�������Jj&#ɦ��xy�qo/�u@���}�2�Z��Xw-��
��~a��ݱ3S����!���8{�Oj1)jͪ}������1�Z��N@~>���Ǎu;��^i�u���k�w�Y�W�V��BI�ϑwU�0��o�;�X˞)j5��2tC�Z��������1�i�t��<zϰ��n̟�i^���=r��"~�*2�ϾC}�t#j�Q6]�VWp�O���Y*.Փ˓k�4V�U� �̊.#�"E[��Ժ�_�MOFO1nd����},�a=">%z��>:�H�m�՜;�W��������h��gM#"�%s�v���A5��Ĥ��yS9R#�+�̳�<W2�L2e|Zb�)&5�7�
��ZQs�o����T������������Ԗ
R�w2�c˟�Ψ����_~"SI�Z�b���|��lpo"�H7�M���������6�" �xB8UVa���3U:W��8N����C;���M�趐��`��B��y����xl+�pP�>}t�D��f;�&0�o�X����p}ӏ��O�ľl��Qy�����Û�;v.Y�)��)Q�k��Ҋ�TR~OJ����Ju�����EO�s$�p�ݠcG�[��:U��S�2�E&�<�� �zgT�A&R�$���!�F���G

���f<���z&��i��G�/�чz�G� V�+�I�?�dnN�#�{�t�J��� uMPo�4-��"��/�������}�v=�ti��w��}"e��5�;zhb��5�c�(D�(l�gy*Ź��Y��LPX��
�d&���uBTg�t�G:�H�;��:t�ۯ�^7!��9s���c��0o�(��t���A��W�8�g�k�Ӟ��̘-%Wd�����c���^%�����	��W�J���C�u���5���W�p�y���4�0��:�#�9������E���f�$���ᳪj�d���6iRՈ,s��<�+���ƅ/� ���A?����������i�Q��[�?6�@�@�s�!�ضq��j�
D'���նM%����<���ƣxnf�������}��x��I)��kr�s+�BT�E�)!��-Y�by��Wc��?&��t�.�L$2V��~N/3 ��9_x{�-���{��+fӒ|l�,&����
v�����=�0�N�x|�|*���������l��#I[nX�o��tG��@���������ٰ���
��M��4�5�O����6EG�xWV�!Qel��f�$���E�񊌅�&���/�Q�+�.��ZR���a�k�m�� �e5��%�*l���fހ|����u)eMJ!է^�ӹ~�ȧ���;oӿyq��}KN��{���8�^7|�!#��<��	�#�tj	*k3n���(S.�Z���O���]2�ЅL���A����j������L�/R;��dE��D�xu�6⧲k��W舓�zwTb0MNZ�O���.Q � ��'M����h{�'��L��p������m�����l��j�'��D�h�|_�cg������r"3��̤��02����^�������!�ol-s]X���Z5�
�1k�|���dv"������9	�$N��.hA�
V��:�\�� ;�{�����á6M�����M2�UT�����y�}oWK���Nď��tX��9B#.]��8�o�WoT����z�	�H�b��
�J)�B�v����j�Ǜ9�������!T8&��(5�e�������5��-�3�# pK�gG�x�)]���Ĳf����	|�7�w�N���
�X���2@w ��A^#C��o�	J%N�@����*X5r�єI���Q�i�T5_zv��0>��ǽ��	�}�7��&*�#j��@�g{��Ϲ��R��x[yy����
��-M�o�s~�`���N�EF�ĘXN� AʝI�m��պ�ⲭ��B�@��)��p�񢻮�+����(�tL4��kF�����p��d�3�#%��Y�p�Ls����-���5%��~K��!��`�g��Sa�� � ��y�ɟ�h���=�F8��J�W_!���~��䑑�"y_��;��rq�.�_T�8�kJS�O�E�K^���]�+���\a�����!6��k?Z��j%7\o�@��E�z�+ 9�1 �N�b:TK����)��Ī�:�O��m�:�n�0�`ޟ�>l�R��:�`j����|ޣq�6%�%�S�0�Pn�-\z^:�U����{����fj(����\Ao'�$ 5s�P1u��rb���]��L���sFfe��w��:a��3ڇ��:�T�7�^�o�8��ЄϛN#S0jN�wlM}�Y�|��F��r�W;�����۞��*;q2 �}���|�!�>{�ɠ��˵-�0���)N(���aj�lBD�&�o)�ɩMK���u�yX[a&�	�T%�R)h`dT[��D�k*��li(�Ё�����^.�ԭL��xDY"���o瑻�?�Rk1Z�'x�]"�(�q�G�#����ze�r�P1�X_�ÿ_t��NT��z�~�������i~�M$���8>�I����H�'Р,���!$ݗ8s :Z�H���ؠ��5�OȒ-MX�/��h���m�䠄�ʁ'��I]��m�Ρ����h��ekHZ@xqɺ �(1Y�S�s�3�a@���ज़���ЕT_*,{Yاl����TR����U�a���E�OH�@������\�q�c�w��q�W��B2��1;��Y Bd3ɤ�v4v+MU���W=���@�wG��#v�1����Z�X[�n��4B�7�"�W6]Ƥ���⥦5JX S~f�K�H���-_e����1�+ීm��aP/:
ѷ}�0}P�q�g�<��D`�W���@����sX�͆q@��J�Bp�O�F�$��L�C�M��U�ӥ��~kN�n�Z��$��AϨ��P�4��.L
q�~��*}�\�q$����(�+/I�o�x��_+hwS�L��0�P�ԍg���۔�ݵf���A��ӹ�'���d���s��,�2��D4
�DHaJt���XS'���R�ZQ�z˄���?!4RɗҋLg ����E�T��K�%�d*�SE?\�O�^��r�?�7I�"@A&UqT����>�}T!�r�?��^[�j~�BZ3��ҋ�;H�WX3qhѶ ��D(#�/���S!edU˵�~
#���$���G���<_�7@PaQ
T�?�2$cݣ�K$��c[�2�~I�'�J��Ԅ�?"�H<Z�����]V����Xw��0c}�d/���jT'���4��f�2���4b�/ںf(�F:����'1��B_Q���1�Ǿ��?�4UEz��w�Q�N�;Zs�l���I��~������R]��|��~�	a�?q%�GQ�a�Ύ	>��j��q�i9̄���=�m�|~���襖w#�i�bU�+4& '�A21��R`d�m�B-�����C���WٮJ�CX��()U^k [��u)k?�÷�7���Ϣm�le�SƓ_�p��+^<�q+	����ΘrO~���;�L���v��Q�?�h;�4�+̴�
��ÿ%�Xj+�V�$WVD�hyq���aQ�y�O�x�R?�Q�>,�^=�/bs{�F&�d����`�	yseev�� Vb�wh	s��z�/�=�\؈��?驁ܤ�����F1�5ݥ��eb-_1��ۓ7���u7G����i2Z���?��Ӈڌs�p	��+���>�*��\�Z��C
��z�@�<��M�qX�����!����(���% � ��6����C�ܿ>+yO���3#䧌3��
�ޅ��+cL��kZ_��T���3F���<�L��j�䬘KLޛ��	CE�P�����Ѱ̕a�q���(0�/�&��Ʊz|ӎC0�u����a�Jl�W��"��r% K�7Fb�`�A��gL\���ny��J�tS�Y���'�`���)��ӛSL�+b�*[Շ�\y:AK�0 �|�23C��]Q���E�3j��tG��̬Ja{� �)T�%>�fDݼ�u�^En�H+̖xp����sr!�����r;�l<吂���<.d��.���{�sA�e��H��F�[�*�j�h0ez���By-�����_�._�����-�DY����j&���v<�u��0�����˗fv�f��[���Lfi��΍��u�A����>t8�C0���jZBE[Why�6\�kR~����⚫�/>۷X��U_[��(ab�pB_!��pwiB�d"�"\�.�#��ʊ��t��xk>���ë�^��Zca�D@����d�w��ڦo��w;{�sòD�6�K v2�m�)���;s�wb����է��a���!:|��?��Q��eaO<?z�b�~W9���z�Z۩� '� �T�0
pqV~IwW���Pz,�v�C}�49b ��Ȟ1�ħjƢ+]���d�L�'>`Ce�8vUr2W�W~A����#��˗��x�.���,����E���qC�E��y%�j�;�}�ˬ�j����\�5�}�wA��	N��)���^�b�lyLu��iG:u�i�)u<�!�&��^ n*�*)�H0U`��U��r��v��Bc�[G}��q����O�z�\��nha`g����q��	�g]���7p�@hG�vR�uI�B�p�%C��?�o�3z	�\��A����g�O�Z���g��Ti/ j!H��y�O�o �-��7������/5�
���ͦ��Z[+p��Xqj�'v��oc2�%����tQ����~Zi�j|,/��%j��-�<m������u�s�ۯ����t�e���߅����]�rQ}F��-y��������{�蘴!C+���E*��騐��$'��V�w������C�?u��o��O�!z7m>P2�E��_`F{�O�Z�d��ݳ�H�Wjj�;��0j����*�*��f͘����Z���o׳(.�OXs�l���M�����ՅAW&- ���I9���g_8A���6�đ�[��l
�釅a��$>Uꕎ'Ä�&r��iq�X�H����y�Lsc3�ŠΔ��sH�"�$�95�_B��d����d�U�G�JS˒ |>�o1\#W��[۞U+�]���:l']����V�(���)��8��2y���������Y�X���D��h���h�+|�W�_� C�wn��/5ȨO���,���#�U&�i����"o^R�$2|��%� aY�o�T��T�1#bێg���3��ײe�8��_�6�n�� ���!�N�Ҝ5��U�$\\�_0��U�:���S�����E=1�3�%RI��.����I �WH�E04D9o��"F�튕!���}�m�%�T�D�{`��1K�+�����Z�Y�}=5�����<����Tu�"���=K�Z <��6�*���JD;>�";/�+�8�NZ�;�F���le���Zx���'�pV]��ow��i�6��%ux~��y
*�-'�_
�3�K&�}5VZ���_~_b��~��ݱ�b���-5^#��>�.�7������{T6#������R22��eI��q[����d<#����[t�8i��7�� m{��B�\���S��O`�=��y ���x���l�"&;Z}fS�ujH�A@%WX6��Lrs�%<�:>��j�W	<�ܤH�rq`�5JkI�Bb�i)�)�p��q<��|u�j�Mg�����7�7��Q�gk�0A�T�WEc��˾XT��&�^r��t�['�*v�(H"�����Ƭx�-]����te7��#�2C���p���;ł�Q���5�/�n�2�
����lx��@p��^�܎q<Þ��'4>/6�T�Y*vHU���'�Ջ���:�pD�Wf]��fQ�H��=4p��#��7O,Q�x�ة�3��f�t�70����T�(t����f5P�2��^dZ$ů�v���L���_�`�i�����ı���~A9�Aȏr��r����q>�B�JXnQ,?�֚qJ�O�Vd���l�=�j��eKaְ��X�4l�U����Xr��^�����}ř?q�
jOS��֦�?��:�\��t��y�G~ū�d���s����Njݡ�l��h������F]T�C ���Ά�g?�X9HD�A�|��+n˛�ڱ����{��ܸ��7[�i��]HX���ϼ�oB[?��=�Г�������X�@���c���׆���R�XK@}�8WJb<����$jd}��v9Z��U,3��ԕ =�C��',�B�6t��"Zo 6�na��+`�������8��~� :�ej(�5���E��^����QM�pj�I���˲��Í����4R:�L8=ؿ�&�x�k�=XW�1Mڧ��9�s9I3
�>}���c�tQ��W$b�;�D4�F���n�IJKi½bv�

�
?�D@'�v�o T��s�;��(��i���hL��j�U�Ҟ�tjO����<	6��!Ɛ�C���,M�`������tj&��zEo>�s�'��
e���J����$}�<�8%�j�ëG
q�&&9�=��wqmv���:��S��	�JFC���$B���+���:F�	�g���K�F��L�#���^'��|\Zw[�BE�"L��K�k��,����<*.�f�j��J���O�	��v7�.���u�ũ�Y)-?Í_M�~��=��[�"��F��Q>}���Q�o��\]tͅ��BױcO�N�|���d""�p��/�qw��01��F�sli�ā�E�ذ<N�g{�7��|���=q�u������0���O�+���a��F����HN*�`F�^��������ѹ�>��G�ݭ�}.f"w���`�D��z��~�j� �oؑ�&�,zo�����|���<�:=��$}a9pqpF��?�0G��S]��lЀ��O~�M�p�x�,�X>]�P�i�<} 
Zͯ^�R���8<6IQ��x�ZՏ�k'v�+./g-]�+����&�5�W���ֵܧ\��^�ء|O^M���%?���>ǭ� �}ωՕ�̖Y뉐�(�syF�QKg��ݯ�JD?�&���q������0r`]�)�,��5ED���)gB^������Է��6*�}U3K��N]�������z��d���RG��ۼ�Z�K�4n!�Җ��i����N�^��T̢������9Q_���wŐ3�;˴�spKB!3�&(BwO�6���*��Da��fq-�o���R�_:��wF���>��?���&(NnNnzSĚ���^q���#ˠ��4��Օ��Y?��4��m��E��j6J�^Ej�r�sƄ�V��E ��%	�\M��n	��'\�e���vp�)_�zW�Ԯ�Z`ez����pWwsu��I|Ye�9߅#�ː����9|���&�k���������z\5��g��<Y(�ǥfN@�G�r������ra�%��s�D������R��rJe�N�_���4p�%{������	�(d�_>U��NA�T&H7BJBlD� �z�'Ye��#��I\�s���W��&��!����gI٠��ai�xn�upA�⧦*�?((�z�`�G?�z�3��Ps��g�#�Sמ�)$��6����n�ۏ���~�9��8���)�{1Yua��3'A���C���"#���Rb�u�)��Z]n�u$�mk'��,��Is퉫E+�7��}�X����"{�:1䵬{���;l@��l����4�~�F�x��i��}��"8�����-��׹qa�ӗ9���@��K(��s5���e�)�e���������Vtt�-~A����	8��Eny�#���I�G1@���}""�e��\�B�w��b~�)��? c�����~����d�"nC�ѝT���і����%qt��e81z�i��I4b���S�95ٯ$>�����2ږkՀ�b,�|J/r�-��U/�f���^��wkkh"�%e6��������`��
k�6�|t�ǦG����6.c$>�V�6�č_�)��i_d���L�mFN����q[�I	�_��A����T:�b�4/JX畯9h��l��g)#m,�"I�%a��I���@c}�k�3��7 0j��i"����cq������0��Sl�W-/��脢q��ʤ�w�,Ш��0Q��\c�tZ0�����5/~��ȼ,���d�����Ƀ��GN�Lyb|gK�c������_w�s%�:���?Ư�� �K6]�ܸ�/�'7�q7�N��o���/���$D��l��v�G��:���c����*G��4���!�8���g�~^�@�1��#��\�&�@�����g�)�4�4���kgM��~!%~�2-m�9�@��.W����X��(	����Gl����~3�u8Z�T.-��	c��Y�	A{��+��b-7��J��{_�;ѫ��$o ��J�@�������v���E�8�߇�Is5H��(k*>(�\�P�؂}Ip�?��l�w������8}q��H���]J=Y_o���:�O挶��Y��ڋ��,��$(�3�]����3�0�w̨E
A����R�&
�����t�ΫSz���$�##���f�Ҕ��[�]��V$ׄ}�������y�0xJ+���&�e����b9�f��tr�[k]ǳT/���
`A��e�I���	z+�����>Av���"U	�~��-�:jkz���G^A���������4�QG �!O�N�6&
�ۄt����T��_��o���	��R�~�^���6�a|엟�����%(*'�X�C�8c���y�L�:���_�d��hWV���2�%���v���z����Sz��%�9H�T����̷��H�-��!�(pYLc��6#�&�hin��K�c�{LR�LJ��F�o�UV�����`P-�����W���^�=����	�?~�/+�n�!���Q%�=3]�א�).V¼���נ�V'��~����(�Cvw��d��x6k)�I ��k:�_�#�&b�,Z�RK�$�H�f������;s�����	���������=���'��;`N;���?�<;�i^ "��# ��M�����&{2���e�_L���[�9fPs�"mo����p�닭L�^�]�`ljR�Q����-f�C�E����9;٨��9PxG����O��eӫb�H�	�:�%���O �æĻ�#��:�9��_]/�E3�	$��������-N�-�DX&F�G��ո��6�X�{�w9<҄n�	PoO�C��o����3n4�1|�1'���P������_7��x��<�`�	���~�|y�4h?��ELEUAF�#7r�yR��ǻ���%��<_��Ձ�W@�m[W�ee��'g-��AL@o�X����P*I�s`z�1K�(���v5#üZ7q)"�>�:I���G}�p��qf�{i`��V��u�LL�򂗼^�LL��(#�*�p���H�o���^�u1���l.���*��*�F�n\�]x0uoa�1A�������ƞ�k��w���l�Z�@*���J���a�]������љ,�*e4u���A���*:ER�Ô/D�^}�>��_,��$0�ᣋn���d�ɓ�M�s��Lb�
L�5���4���9d	S[�(:���h~���>��/9,��%q���;��s�\Y����JN&S�� T>�,�Y��)��h����=M	(���U�N�Tq�S�r�9��8� w������.�:�A�wy�S}'u��Ì�`=�����@|Vp�jH�e�����{��v��Y�t�ɓ9�c�Jl4��*=����J�}5���'&����� �*U�*��=����>&�&���$&�?�LF��,ݛA�>�.E�)!�B�]uE.`G{�qZ����x^u_sM"��/xnY����R'b��*�_��!��x|I�R����q,���|�Y@f!�:�����[+��V�t��{E�̴ȣJ*�D+�������@�p'r�Ys�q}�O9���S�Ԗ)l3_�C��U?I��*xӁL���ʓ�<�O����;��7� Q[��tY{-v���`���+��?�J18@Sө�[P��������?��Yo�����^M���z�>V�	���X�gcPT���L5sI���+S�B>u�0�c���Ў%GRf��,\z���WՈO�Ah|��,�Xr2���n�I�65	�(.��d����E�5�a�}�����*�\^w��jd�}���	�Rj���P9��V�u�A��2��o(VS��u���n�B��=У��i<�0+'�zWI��y�NQ�%uzA6�bƝ��wKO�o�v}�Wl�@��#�����IyS��d��r�#Σ?f
�bO�1��Y��%l���)I���-��S唳�d}�E��<*�����obr��nx�n��QdL�U%O�_�-v\�҃�^jk�z�A�;���g=���~��m�a²����SwcPس��Ŗ冯�/�t����8�۲�**�gL�$��(�����<#�;
JvD��S���=�5�TPl����2�:DZ	���>����ȌZ�)|�v<�쓔Ω��&z���rB�����( �R�/yqP]�2�ѵ<���$�IS���K$���Mc�샴��5G}N�ͪdd�ʓF�[ sО�2���U[��}?G��k�;>b9>]<�J�����+�c�`P�Q>�B�KXg*[���1s:A�$�)���U��jBW#ϋp?��}�a�%��*����.71a����E�r�dCum��]�⻳�y"��j#��$���-^�� a�U����v��sV�= �o�ڐ���>X+�跠�I_o������¹���H�禪J����S�I��"����Έu�
w������a0�B�S\�r��m���t���Z��CS9L�k��� ��$��X�j���!Ͽ�Q��;8o��R���8	�54��_Kc1P2�e����$jߓ�KJ���a�����R�K��Pz�k�`��z�7���޲/���/E8�F�[�=��� W��$bKg��H��h���4�=�ⷛv�+Q����2yώ4���d�v�� P*�c�Z�Ƥn�����g�5ٵBd���@�p�T`����\#�3������n��Wf.�@yqAɰ�\�~eiM��D�&��܂���'F|<,����K��	� ��_�
!�&�N��g�e����촙��(�bt�']�Ր���d�5�e��������x���0�̦�բ�x�}�~�>���������Ϝ�&��"QO<���d��Sp�`�@g��&������xמx�v��=%y@��3�ۂ�'�0h��v|�<D5�Ö�wi��t��l�%i�"�_j)�ʗ��^�܎�?V�`Y���G��U�D#szo Q���2
OKۄ4BUu��/x�1��|3�'�<8=��*��W%ɭd#d�:�����9���D�qA��}�(D���P]��9�Kb����P��)�T���B�����;����ɐ���!�����	��~,2�\��Hn9�D�� Ҝ�_�UJPyK��~F��|�	D�J*��9���.��(�����h�uƨ�
N3��d~"��mC�����)�w��+��!h\��nd��y���-1��*�9��T�����;��ax�V���ww����R/,���/} ������y-2��zN��Sk����B�ķ���<�۾��Å�M�[Zc�G+�w3�̈ܖc78\�J�w�s�"�>
�-$j�X��{��*���ELɠ<kq��|]����G�+z�p��f�QbT�p���5��!�>O�������}����m\�J��B�'-"9�p�/S?X��N��xO���4
u�}"u;��}n��@��2M�Vü�2���z�� φfFh�y����-4�V^=;>�X��_��x-�:�4���r���l_@pI��a]�?��A]
sl{� �?�F/y(��Xw ;�x~H]�'�4V��x]� \�/����ycs���V�X����(��_�jm��	1��<�����vB���ŒS�Gi�E���g�Fɽ�ǰ�45����7��a}'�7�C���`�!)R��g�8j�̈́i�������o2}S���p���3
��*(��}W@G��1���փ��(��T�u� ��!���Pu���a�h6��Y6Od����%�o��P��8
�Au�� 
�g���	��Q� 3�1��O-����G��������+�,��׭;���_w���P�@#_b�݊k
�Wb5��dTP�02itR���e��%���6�fe���8]EՊ����IEڠ�p�w+C��9{��܇�#�<��l'��<_��{��K�>����X#����0�w7q$������dc�>��� 2
�4�;��́6��T��5�.��gE��k�W�^'���6T^L��X�)���L_*�M��M��O1�v����%�m�?��,,�+X.'�-~�9k�%>2H?j;��I���o����c6��~sz2C}|�k�UQ֦6��h��_<���^��>�q���\�Kn������yŵE� �_L�F����Hp����
�#��t,p-�%7�ݾE5���D����T_~{�m�$[�j�`!���^;O�_h��,jji�澲)�.Zz�����4������k���,����N����ު�/��u8uj�^�Vת�=k�P\Y��l^Y�KgLE��S����/r�~��Byʗ�K��h"xTx�= ������[JZ�=��yA�����=�M���%Y�o���M1��_];a��(��*�*�3iHǀ��+����L��?E��bբ���m���h�Q��D��x?O��Dĝ�=C��qW(�G��o�懨�̫��w�y���7�Y���va��#.���~Pq�!|bacFi�Y��+�$pk�X[�����<ݒ��J�����x�5�-���JT�^����::�@_��/�R��--s��s�Ɍ������9��r�G�v���]�!�:�<��M[H���3�� �u�2|�[ʂTS�䈖���@o��XV�<���[��G<���ؿ(�nSݞ���K�@�?o��V�/f<��S��g_n�@�y�f����Y�9^���e�t�%��{�I�\��u!?�s�[V.�K�??����=x�
�O.�_��1=pG�mm,DN�����h��h�X[Ý�e��Аd��$�2�NQ��~���&��3��{fG@x�hJ���zh���.b:5����V�63qq��W�X5�i���>����I'ÿ��ټt�/�P.º�>٧�8Fɼ]�7��ζ�LL�B� �	g/�S�͡��rZ���_r��r�>�ߊ��8O�L���ر⓻9�>���PV�%�����O�K����JO/�dP��+�w���A
���
��yH�O&�t��T������;�����V��G�9��LAu���w�i!꣱?}���;���W�./mą�bq��"C_�Z6?)PS�u$�P��	_����Jk�ٸ�K (U����A����bu�O�0�"�JwɇGQ�7g3� ٷ7��C1�y�:(�4�ȷ��O��2	�cq�4t����ÞOJ
��0�B�9|�W�/��D�ە���,�#ֳ�4(�����d�Oïе�fb� Z�%&�;��pv5b~df��K����XrV�+bc*�@�ꢂoJ���&A���@1�o�l]�~�:�hyY�H2؜o�r�&=t�s7c�uQ�����p_Ԩ�D˭Q]�~F �o��7i�����|�^X��>U|�$�}X��-}D���C���J8\W����iYW|����9���A�ֿ�����¤S\�e� ���q�:g{���Pv�"�+��G�!�����^���j�@�	.a%F�g��Y�_!�E�q�3��}<�����%��ӧ�hio��3��J�<��Z1��b0�n���%7�cP�Lb��7.G�8�Ѵԭ(w��}�ޙ��=0`��Xvl�%ɋ�"�� �P��n��L�!G�Ȟݓ�IX��\�`&�=�g�-AN8&/��ya��֖�nއ����Z�O�~��x���DdWߧ�7 �)M��0�Wdh�����j�/BH���e8�P���p����x� �Q���-�|,��b�<@�;�	�]s�>L��t܈�a�d�K�m��U�CE6-]$�:ĭ��}��5��r�]�e�Ab���8�
�ӹ�>�1rR��g��I]�J���_��O��+��юg�Ƿ�h}?Cb�{�<���a��M�3�O����|���y�_(p�,n#��v��P^S~�����Ot�]媺�B�Ʒ����w&�u3ѰDS@Y4(�(˵#/�\Xgu�33��s���x�,� ��n�m�A\�h�1J8�%,����D�Z�CR�}� �>�籀�y����T�>�g���u�^k��ASl��,�Bĸ����H����/LBb䷶l���sX��o�2�j�_�ߖ�>�nb�J*_����\P1��)$�K��R����+�r%ުK����rz�mf���(Uo^z�_=���k��k�����M�I�� �lT���� �X�g����[w���<��z��!��V�{|?w�߅���g6����ۜ��� |�.lk�E��*aOl�,z��<ce�\��,yɧ;��"�ڂ�Oo�7]m"Vv8{����0{/��A��D�F#������vm1G�(�L�j ����xϩ���F	s�>���-�Ls���Z @+�fL�5��^���J*����)�1J/<�?|�	���LP��b�����w/?�p�0��0��e��W��E��H��u8E-x��	Q!J)���z�n�D@[1��5�P74j[�:�*�ڝ�*W�~E`�gw!��1���!^�{�$���kl`�5@�yv����3�y�_9���^bVĿg;"kKǮDf�D�!&�.]~�F����FNpa��m���xܰ��'�!hl����]�U��Ⴓr�]�q��<k~֟�{89F����U,�(Gs`���b%�=�l�-���1[�JW¼uB+�O�2��N	��u�J�1��g|�	��>�͙�yi�BHu:h,���]*&!-������ ح���!2C�<��e��-¾.^�ӻ�b�������_>�@�j�qa�S��o�����R��p�o !%w01ܢǽ�D)h�V�Yg��o�;Tp)+r,���b��b1��/�gF��Y�xU>xnh��� ���Q����a������@a��|��N��� Sm�!nF"$��o����+���:�la���6��Q&�w}���F}U�cTuM���$`E�.\�cd�!�����aM��6�k�VׇK�����P�
F�؅�i��� �7@8�/�����h�G���}�WE9 -���>KQzkj���/�P�G�N�!�{=�y��W��k�!�Ԋk� �"���V1����$:$�CZ�a*w�.w��S��5�WYO�٠ZT�WV��U��P�.<����5��q��X�qIw��ʐ�B�ҷZ����X�R!B<^�8�,�}�Ӈ M��i7������
�\��ԽB�Ρ��Ϯ����x٩1b�dX�ZS�_�d1�-wm8��X�Ѕg�@�nX�A�������W��͉�ee�m���f��p��ZF�-����2䛻A�*%��Cy�vS�~:/o�~k,;�a�j�L�	qf�Mp�4����k��� �����Q�Y��h��)<vŢ�vr�G���;�g��ٜ���6�]��+��^���N�5U���-�g����t�zbt�όq�m�7wؓK7�ᜥцC���K6�!|������ٲe��b�0|]I!J�?�V���9[hСӜ3����:hS9/!y���h� ���byH���w'֍���4^Pg.�{�8��E�Ҳ���8�n�"��+R3�]��������m��R��n	�Z���E�%۪ XB�=�Ilj=�trP)�*��9��2�(]A`�� ����Wl�Kq�_j���,/ta"�u�W
c91tEY=Vk�:����6�ޤ@�˭��0[�ћf�Ǭ��=���N�F%~�X�E4i[�s^���-���J1�oy�e(Ek����3�i�;0��h�%u�J7J��y���ڶ�o��\�263���o���|A��ҳ\�c�D���,l'���ͷM&n�������fɊ�f���EXʪ�̊����Z4����C�I�EBÌ��m�	���,(Q���&t`_�mA���aͻ���B�M�гb�8�Vq���,ȗ���L�W*>�ޡ}uG�ʩ)��)U�޵b+kT6�}�S7Y�!�{"�jǏW=(�}��)6t{��(cz+��i�����r��E��;_D7n)�}-?�#�̦B5*~�W���}�7�*�Rr��
�Ft�lT4?_5b���/):hB[aJ?s�����!�������]�:G���6K`���8>!�
���m%�Jޱ'��}����)��B�X�J��ƥu|���|�:e�ϗ��n*}��?�6���j0��Ղ�d���h�Vk����ܟ�_�=����_�Yx�XQl`v*���x4.�P���R,��X�1@�>����]���G2�dt0US��\�c/sKU��X�yG�V�($-��<�{&���d%^P�ńt;�I`ו�&�ύS�*�Lʳ���V)��[�\�~�B�2��}%N��#!!Ռ{��cT�8w0�֖������A������E��@�4�����~Z�/񝩟½��}�R%��)��*BqQ�����K�FJ��ɋ�$]��6�W��v�K���Gwb������LZ���F�'�g�Z��<�j�6H�LdBm���*���Rñ�Nx��Mr��Lc�^9ŧ����>J�껽`��w���
o 1�G��m�Y������9�������|���m���9~�W"�N��������7@dQ^b�@�,d��M�� �F���.������d��K��mW}*�#�-���8���`��$6��s^aWFo[h�	V�B�	��+^�=A�;��a�F��A�OC��\M����g�O�]骄hu�9�����|���og��]@��j��W�\:���J�L�ϕs��Y�)B�:l�1�L�vT�%��T(�������$�sc ��J���N�RŒ�I�*�H�J>���R���I��sZ�ď&_=,hn��Q#i�!Z�z^������}����9!��1G÷sݒH���m�������wt�}x=�����,�i�z����s9�Rw܍μ��^W��2_U�>��S;��G26�8݉rϑ����h���Eq��|����v4�.g;�.��G��p ��{�;9W�T��/?��� 5�f��vf��U��_P�_�x�$�C��:>hVL
�T�)����h�@<`�ww��e��ڈ"K��f�AҀ����a�`��,� ܟ������� 3�N�&<�M�K�5۟L��c�MX��c�^��\�U5�_����q^��%��7;,���LKp�[�^��K�}d1��ä�ZZF��+� ��
xD��������	�w�[���ҊgH���?)�?�zhI��u�k(���>��N ��8�I=MS�<�+'���8��U����FWO����:@�\+P�28Ӗ��`��$�7"2���x\�
�W,<�g��X!��->=�<�Oq:`����F�p��ar����'�Q0>'��K5	���-h��*��Ƴ|B��ڟ!�SK�e����De4� �~-�:?k������pH��W>��[���*�"g�޸ �T:����	y���7���w�Ll��f\�f��^W&�x}8p�R�l��1hW�og����*�E�rM���������guXR����ی��4��%��:ikZ�l�GQ'r�ş *�Ƅ���x�z�ݔ�V�Z_�.o�d���}���Y�;i���i�4gJ���K)yQ���1�Ն����&yV�s]�����`̱�t������m!!7�� �.tƱ�Lx��8����T���Oӛ�6B�#H.��z��VbO�-�N��4�t����uI`2�JV������N�QC�Y�VBHd���D�$�GR~>`?"h�����yz/(���>T�&�:�k�f{7>?�[>x�]lP\{L����Y��j�9�_�������0��/����"�A�.j�`BD������xz��A�h��o.�����&߈���V�}[l*��)FC�H��̄�p���F��f�� ��b�̀0�k��߄߳�u��+�B�G�~
��=�?^�[��PM�6$L��'�`����YVm_���/B�A������K?�ɵ0���.����n�9�
qqi5|`A��՞8X����O�9)5V-��Pb���H/�%Ln�vB�X�x�,�^����z�\���H��q#� ����y4�"%e���$�*ǗJ�0���F�=�u#xt���R"�� ���*z�x*���~����jb6pЍPϮ�zw�mѬD�WS��Y0��I���祓�w���z[�dK20a��[^*�e�/7c���i�w�X�^����f���!0F���&xa�85�6��K��wSR�ǻ��߂��%/t�R{�%8�d�U���w*��6��fA�6!�����5@p��<�/�%G�;F?"��xN8�8����PO��s��-����mXA2n�N|m�(W<�����"�i����o �g�#D���g5�}}�n4���㧧z�o��r�|��y��:�ge��&�K?D�,�6�����⩰��?��5	X�	�'��=�ȇ�J�9��P�NP�>�d�`���H>đ�	-�(sF�K�St��mG�i�'���)���Rfj��L�q�	�ff<on�0[N��')2H>2U�~��b����h>
�W���h�f��@_0�%hzq�ۿ�{��~X���
�1�;�0a�x�>D�j�������t��9�x#9�boX��xH�`�*�I�E���ax��=� ��7q����lpؚHЀYsE�,w�=%6�FM<����j�{�x��>�v���mf]Qf�R�"�o!����̓�*�*=��A��e�*��m��jvr�;�n�.���N�F͆*=2e������wT�녭��z�%��1�J1!��G����6�/m�X1F��F�/�`�:O��@4�d�ASU��r�E#P�B}逅�|e����γD��*]`x鵕�e��}��ŉ7x�9� �
3��I�q��`3>��E����r�O{@��\�<y����g���_}���]������+j��[W!#��BÂS<6@J���8C��u�X����'�}{{������;��t��z:3�&��.J��K�S�$�F9�1Q@8ﯔ�P�ה�
!5jpZ`kz^m���>D���y>����ֿo�0|"5��z���Ԗ:��9��+iU����[X1��Kݺpv<��
��M���Vަ��pr)^��!�T��bB��2f9)W�B=?A�c���yjof���ֻ r>hqtI�p��ɉ�I��gZ�]Zv~ʧ�������rԕ�ˏQ#c~ ��1������r�ʟ3!7"6�,~�Ϳ��l�1WM�&�	0��
�q�΃Ǳu1��L�z��z�<H�*�/j��d�b�|�)��3i�s�ՎO/����E3/��C��vN�_�戳h7v����c$x�u����aB������z�u>��V���%yՌ8�ն�N�-(�!&B��y,d��K 5y�
?z���0�g,�^����0��k�k��D���Έ�7�ɺ�.��(�ˋ�})�	D�t��r{��Q��\%6J��I� ��Q�0p�4�x}��_)�0ӓ��L��4_@~a:�9�q19�ɶWR>����N) �	AP{2�����D��_S1cC]ֺ�c��_��^|9��u��	_D��o4�j�� ����x����������!"F�陵��l��FD���;Wi�*���#�K�wzO3o���1��^��q$�����Ȍ zG�P�0&�(R��'�h_�Ƨ����$�,�1��ZO�/݄�c��I�4�/#�����o��<J�$��-�SZ��V�'���d��h[�Mw[qqݰ�!P ����d�7��F�E��׶��X;�w��*�)��x&�rOh ۻn���[�t�vV�Z��V�e��ه��p�J�p�j�f��W�'��u�8훁3�?�L:��e-�#�T8_����vg�� Z�(|~�(r�-R�Ǹ>K�U�����`��9���t53��-cZt&9T*��=��}a�Μ�Y��������"���b���������F�o�����	6P{��K�����h$W�T��<3�o�ܰ�+���a�泿ΓLyYQ�G���v�}Qz��ur�����c4n@&�D�'R�0���q��_j�V��{���;�s�������nv�im��ş/�K��q�^/k�����S��!���C��r�s��T��d��w�y�D_z�D,�2g1XKQ �R�l�S�$H[�J�5`��殢�.�
�m�EN�!��Ub��EK�8��$"t��O�ɮN LGt-Rʡ����)J�̨��̫_έ��*��+&��s�w�1庇�y�gg�=�XZU�:G�+�
D0���Ʌ�&�JS�D����t�(Xo`����uw�)5*#���X^P!�P������9�KNZ�x+���۵�/�>�_3P8��P]�7���H�[�3"P^^J��P��D����j_{�Y��H��e��<?TkH6xpު��5�frhjV~g�w��s�&�vf� �-ފ�U�(�l���A��ܷ�?���d��(<�˂�J�:�-*,'_�߀Od��Jp޵St���4�� Kt�5y-
����l�VѠ30hb���Pht�Q;@�3$����rP�i�.��"�|��z����F�Կz��W��`B�_��I)��d��i�8�MC�o银�+u���`�A���K!m��|���g�_��%�Ťx�5��8�4Bj�S0��?�`Y�e4$G��6B�z����8�쨂?#�������"�$n+�cR��O9s\t'%*L�/ ���|m}��#�ؘrj4V%T��E8
�x��ﵫ��	G�[w�2��Q�+�����q֐8Q�� ���UQ��g
�'��C��$�X	�����r�R�9d�>�gu��5㸸�;ϓ�͒B��m@��jx�HֿD��Q�l*��o�IhL&R�n>:���`$h\p&3�(���wv�{�ioki���� *�9\��nN|V�u4�U��WR��}�Y`}h:0q��O�b����Y[a�jn�h���(�"�K<��7�f���}1{:�k���k�p�nNd
�ME�F��@�@�2Qx��<9����3̻�	*�r���H����}2z/m:���픭c��Y��ek��d�LNK��9L5��?�_7�P:^R?�r���RLlC5Ջ4-��±�x?������_1a�F[����h ��e�'���@�Bu&�7���ӽ����:�Q�2�L�����:â��w�����BP�fv =�s�Pm�V�ͭ��*+�|�ۤ�$�� N��1Ӣ�1u:���r�[^�⩨F��o��ϸ<����i�i{$G1��K(D��U�lF�!�g�{l+��U��f�ʪ }�@�
wa57
���/��d��#���4.����˗f���m�d��J��L�9�9K��T�2�0�R�|_Ɔ~���h���o�b�	�b�e�+�V� �3���u�4���.ÏE�?�E?-h�h�Z��8X��c�
�j�Ģ[���6�R����N��Q��PZ=�}}����e�4V��*�1�h�Za'�����W��~���N��]��ԅ#b������셑�Ox71�1vx*��QY������_\\��4k>��BG� ��uè���4��Ig/B�΄��NXZ�V��2��>�5Юp7�1 ���$��|lk�!�H�%��C�����0�y�b|T��bO\�>�<A,��g�Muٌ�b2�X�.��	>�a�_r�7�r���w@�ݫ@�A� ��<A"Q�ɣ�=��%���%\�c�#:`Ls�t�\��X�۝��ݼI:���
���g
:a<z=����x�,��
)�Ǫ[|c��Vi�l�>4��[�tpq`��rG>�(��ܷ�,y���r>kC�l2d��hk}��Bg x/j��G;�]h�m�Vn��څp�am�T(��^:��Q�.4w ���QA#���q� �U;9�*�\�;^-�w���i����\��۷(C5|N����1]i�y�4�\,�ʐG�<��A�[���"��j��"�<�w}�8�k�*k ��@_��`���/�a!�@n"՗/h���*,��Sȏ���olQ�����(�U{�Ub�G���
Fճ��9z
�Y��� ���m���5,/�:it�HE�`��x�Έ��-E\���L�hb=$�jdH���Fv�H_�(�hk�H2{�
��h��E����8��Z+!�������WM��A�U\ gb2&�+3x��g6�/1h\{D�ڥ����\��SyS����W��)	M�ĕq��D?��V��<f�]7���?��x�%��N��~�~8!3�lb�_�����أ�@���B��Ό�[�<�ZiF�*q?��Y�+-�c��G��U��+��'�'-��&()0fa���A�h��o���O�RT����� G�'� �ź�6Ku=^6J�$��R[����˜wI�@7��և�� |���7�[�v��P81{Q3��˥��e2�5`"��rZ�FChY�B�7��0�|Ri��&�<�q��=�Qw	#�G�����[Q�k��n��7��#e�o�d��=������F-��j����M���j.���4G�e�w9��w7�)sū��?�[?����L�z�Y�?��Q�h����WL)\��7\	�x�1���TE���E�зé�k�ſGY�yQrz,�A1d�����oȼ ׯ~%b^0\�y�\�&�&�2r��aa��R���*QjxbO�{�����(n�}Au�w)��C��<�) �88q���L�.)����P|��*ˢ�2E��دp0�n�Tf��/�Ɗ�z'��L��.��,����r��8=�6��1��g���	MD�������١��1�c�1ꞯ��ۆ�k���n�A�=%{�j�&ƣ_<�G5����J�M��z�!���v򈧆z��$SR��Y�B�M�3���R��(��,g41җ��4�� Q��3��,(���� �Qw')$r,�"h���
o�.��NQrs�*���L�:�zD�8*\0r�fc<�[.�@ʮ�\���&8�:�2w7�ur(������y,� v�����E������.-�_��5^> zZ�	�;�F��C�:Oj�0v�h �@%� �ݠ��=&.΃��%~��������'��.h�U�MA�~��p�`��&�ݎ�L�f#Lg1��Q��ր�]7�Q9d"��S4N���D��Qas���V�,bRL5��~FK�/����j�w���c��ͺ�KDV�
��$�O��/�R�#4�iU��Ю��H��B+��ײ���/��$�G�a��'�+�������l"Z��xY�g����T�z��-�w����*�ǲ'E���h2nԡ�X��>�"L�pi��6B��;�J�tq��A	��n=1\d�&��6cп/�3�؅g��.�cY��պ'uN�h����� �$%^wK/<�(�D~�Ѯ��J�4��1����?�mM&��aN���A�(�_i{Y&��C=�a��E%;˾.�h�>푙@Z���7���^��T�S..���W�Z<	]G�?a+X�='x3�tv
@�R&��꒜f��^�t�Z#)n텟!0��������9����A���������t���^�`Hs��k����D�?zh״��%x	E��1�E����4Q���#��?��2�� rҥ2�Ӵ��N��_�D�b�;"���B6���0� tf�\� I��heS�P]�)i��v���u�T}8�"�!�[�W�DܤӺ������p\�~���*D�*uO���=�t:o�M\�/�i�g�[}�>{UG����S�a5�U��)Ҥ�7�Bڛ]C�0�t�q,Mh�D�ɷ���͋tHLPw��GD?�'�(���j�tO��]�a��O`Wek$���X��3zۨ�_����HC[C�kY>Ek�wC���m��Xh�F�-��f����-����Vn� z���24m���ܳ7�J�\��S�|�$vX;О�*@ʟB�/�?�|GiKT���~�#<��ȁ��J����I�T��m��2���(/R��
Bk��`k�[�^;�5�O���.�.��&y�ppZ�<��=��nu^k)1����W�[����ª?�:ˮME�jO�3_���8��z�ɼ�+߾���?�׆���}�]����c��J�3�=�|sEbr����ȽQ�F���My���e���,�oZLYS�J�%���ئ�ňM�:�>��o�M����0���g���c}v��y�����Sաe��Ƨ!c`�*��������Wb��d)�Vf>՗�C��Y�Rj͌����%T�N������򓆙�N��� ���@yj�,�ZW�7@���;-��3�D&�ԑ���p�ݸ.%^c�N�Rbd��5�x�loMU~�.ݟ�t�2��f�|�x���l(�����-v�VW�����^�n�l�-�hmY�([�w۰X^1<ү^	z�K��?a�{�^����O�����$���v�gP�*	j��H��zVZ:+��L�8�Z\���b��ޮ��7��o��Tұ��}δ�33�>��������:���+39�who��!$�$���:�U?�P�*+�?��x�Ti�p�.��Fڍ����XYHVN�&��<X��F��j�!�h(��d�*�-���#�K��h�'ԯEh�4I9�����w��dQRrT�I.�,�\;��ӧ���6tz.�'����d8/�u�l��+� �+O�+�"���� ���g�6�Ų"G.G�R�L�WD&�Κ4��s)�-`�rztR#��d�
T�Rv#��W��NN5�Ne ��d���W�NG2
�@�:Y�Ґ���M���jX}Q��R�M�1%�5%����ZӘ%1߉[Q=����vb�l���X�� z���R���OבOi���}ż�/?�P�DJSkJ���'��s��Yd�؟���b4d��%#��B~���4����C���ZI'RM:���jxܺ���V�� u&�,�gV��S���S�FÛ"uFJ�I�a�k��K��2�W��d�>�luIx��d�Zk��V������l�C)�5�է�����2�ᩱ� (�tx��1l�9֊��r	"�.�'����)J�Ha�z-{!��Ur!�\��a��a�xͤEy��cZ@3W��!?�e��q��Ն���K�C5S�G`���Ԡ��j>�A�v�A�
����?�����m���#	PG��c�
S�c~���Լ<�]a4.u��W�ƚ�T�y���|��s�%�3S��a�i���F�6vZ��q�N�vy&R��Q_d@M��r����D4J��:�T�ryvK�E8�}�=V�9��3�<�ޗ�@��tb\��I��Ή�WԆ�n��~���kEԌ�-�)ܔ�D���'-�#�����5-�*&���8]�� ���۴�a�NIf��5���?��	�Z:�_�L҈�&3�5?>X�8���/D�G��Y�PMJ��OR�LzN�_�|����T���\f�e+J���^�^4�B���]���4b�t:��s(��>�j��=�9�}���C�K��9�z����2����6��n��7�*E%�^���?=^�ȰQH�\��I7�}�Y���-j�����{=ƇG�0��&����������-���E[���;x7)= L����#|�ă���l��/;8�� 1��
Q���h�A�"Э~0Jgs|pΞ]T��#~7�n5�*�'�Pi)��^*�����������q)!��S����r�SY[����x��:�]�zf/x�c_¦�Ӌ���R?�����a*U�G��;"q�]ڷM�5�06x�\(�)t)��C���9�Z	'�M+�V�W���ӯ
"��ZR�ល'�h�m���?�_�}�֊�[q9Z�?� Ϝ2��q/d~�s��m��t���=����B�b��Pn�CF�e���n���K�Ȼ�-�����D�W�=/pKw���@� ;��(--��7H�d�jk�wQ�j���7o�f��|��8�t0�ؿ���.8?-�����Ps��@����Q
ٵ�Wo��@(���qy�?ز�� ]��'���)��wS�0o���
r��s酟�h_p�?��v0���6��|���4[�c���O� b2�rtW9��ֹ��"e�U��$���>�mtW�7��mJhT,,M�}c�6���m�u����275�/�NG����U5Ւpu����E����OC���b�z�N��2��6Z=�b�~�q�M�K�
(T���{&跎5m홤:lz����y����%�zPY�5�5�nN%�~P6�o�*n��sy!�%���џ�Lݑ����J��a:Y�݀	 K��;��)7�{���),(�g�����x[�.��z8��w�FV�w����~�Ç4���D���"���o�[�H���XҒd��4W���u�&^P�5?�h9+� �W�����"	:�&�5�oW���[.*��ql�Q��i��!�f(���Ԛٟ�q�E �U����`Oe���������%��*��ē$4�	nF���1V8���:~�ez���a������Z}H�sM�V���������?�î`��(�ؐ��>DNA�"�#ɓ��8"'R
]�霉�֕��1@�-?��F��}�;��B%��5^�o��S���#��>K���هR��#N����9�%ͭZZN������ey�BY��.|K�f��N�Ş]�j��0����"r;�,�ǟ����!����sÎ5捐X|)�'����b|%5n 
؆�O�1�S���xv?�VH�)��hmV졮qǦ�6�yy}��M�
�ULo�&����,�[���s���U��v塎���m���*o՗������>)^��
� ��䠁eA�iQ�՝Xf�)!D-#�=S5�����6{����!�$3�Ђ��L�{0�*����IǍ���^rW6ÓG;����P%h�=���P0{_�6� "��1�2��j-�)s��JW��S�r$��
�}�3�5�8蝊����~LwS"�QdcI`�}���|�8R����t���,h�yb~:�6�J6��^	i\J
[WV,��fJX��MN[t��q�\���CGU�1���_�r-��'i�y��6���0~��%ܜ,C1��`A���R�YIOf��
����0�o ?�t���
�������r����B'�n	�燐⋩r�Gkk�a�`>��7��г�C��E������t2���w았=��q���Xն��c�5�	�w�r�S.kׁ&�^����2C����Oy:,C���] �L{ؖ�]��[$uf��֌�M榕��3����W'�ɦ�J���Zх���-�Ҁ{��8%��7�����ŏ�jQ�J�/5?�u�T����7�'x�d�:,�@�\4��NV�A�Ow�W��g�
��y���~�w�HW�m([W�������Oǅ���߹
�x�b�4e�<��
�.��x�����k�4#m GHC��Ud�ۡ2f���<�������_/���
"�g��˘1E|���{�	`�f����FRb�(E��mM�1ci�R=W��vѝ�S�겇��k��� �g�KNk�.�MPrF�'b� P����ʮZT�\�%-el'N�p�]��8RXq����i��/l�������7@d�������Gf�$�e�{.Uu9P�p��AnзGyY&�������ID:����^]Z�?�ވO^;�_v��b	aP}�� !�Q0cZ
�"���b>
}=�b��5`�'��@-�:!E�IZI	��Y	'�:e���z�I�>���0^Ǔu�v����k�b����1��v��Q��iiY�����gk�I+� ��F��&��(S8p��d�FBOԢO6;2��-TK~����ʹf3��ׁ&��k�WZ�%�-#)��Ʉ��
�><���]-J�^��!$��5h�q��b���N�YN�=�;8�<�2���6|�˞�j�Rb.���;�wf*o���$w?WCd����	�����G5�^�#���iYq��5�8l7�~�m�u�!*/�ը�$��]�[�"ۀdT��Z�r�:�!�;����u.nǢqx8w?>�i�L�!J^m�]� ��e$�i( �
� �>3�b̢D��D�Ѵ"l��g�ܖՕ�:��S�&V���G+V^�7�4�Q�^��~����y�ֶi�Da~�[�_�N�/D^������ˋR(�CϢ�K��'��j��BFY9>�X%�">�X!����!����*1�K���sj;�Uve��
pO��p����p��=N�mޭ�^+�����֧�Uq���G�L��~�59#y^W�����J��%j��@ ,�cVVus��qU`�Lv;W�G8�����ܧ�5�RQ��
��EF��Wι]ܫ]��s2���P�&��~%^���?̝eW\M���4��;����=X�����www���4�����;b�{}�g�s��WU�:E�*!�t�:�L~�NN�] �&�K�]jb����
�z�r	%>�=5���~5YBF����	֩�ʷ��O�~��Ҫ20%a05���*���7��4�۟���O��s����&2�~֤ޚ�?j0��
�vl�ޗ�{c�{�s!I�܌�m�G��%�{�ZA�W����Tzn>�r����1��̀4x� ����(��[���� 
5?�u���{<�.���&��1!k�ٽ�n��t�*>2��ŭ�o>c��c��UJV�j��=Qr��Nn>�N�8gMe�F{[Rk�N�ICmC����<NNܰ�4;:2�`�\����YR���>]�ɫ�O[�KMH"T��0�Ě�6�6�&(TVVX�U���&�[�0f���O�����wO ��B|@������\x����=��q���\���Kl l<C�t�8MBN$��qdl6�P�E��#���Cy5�,S�>J�4��~p;&Q��5�չ!��nT�)�	�Y5��A��K��m2q�Y"��¿�����H���Y�47��q���;�0�p}Pa {+"
�����"z���^G����E?�GiQ�zL$�>nB��th�he��,+�v�a�\9э��Ɓ�}�2�Ou�u6�_����h���F��XX�ֳ����'�����"^���ZZ��AHT%$�����͌��9~�K]�Y$6K��.e�G��~0=�&���� }���$~�x���	��&�;]�b]I�Z�h���Ze:O��{�@���I/_S�a���%pi �5"�������=��y���y�x�Uhz�#[�g�=�F����F�T��Qj���!�^�k�ʂ��n�w 3K7>=���;7o28����-��>�x�j���l�?1_.�����
^�-�)�ds?�� k#1R~������YE�VQU�S�E���({}�a��R��՞u?0x������޺��c����=�Õg��zI:kM�ŝ͢�*��|\���w�J���I�.>S���$g
0�����H2��f���1A��ՠ�^���@��ŃĨs�4()���	+<"-�6�Ʈ���nyoa��2xwhQ�����^���ö���$�2?�|�Oy�
6���33��H�6�T����1������c�M�V0��k1QY�ܲ��ﳘ/Ӧ���G��f����-�x~m@��oMZj5~U=I��'�{x5�:���x��"v��Ɠ�����S�%�N8W�"Yp�gd-�x�s@9�>7w>_>J(ے�ْ�E2|��e�i��/N���l�R�^O���2���G`-wW�km(���-������a���H��F���`��h�m����nxed��$9�tB�n[zT�4�VL��s����H̆*H��O) �+!�+?�j��)2�Yq +�A�Aof@��^֝�rOcȍ���y�D"xtޣ�������vg�h��%S�T�\ܽ;t�{v�c�x$�1�(|*�af�\'���#��!�/̗��q�3a�=�s��ݽ�G*	y9�>��E�(e:λ4���j��|�{�ݝݣ��֜HR�)�N h_~��z�!�g�~����!���xH��ޒ��a�b���Y ��:�f�E���#����@��w��X��>���B�|I���Y$i���a��3�j�|��P����櫃���g䎟����ăh/ȷ�j[zd/����g�s����܄I3\}����ҵF�:73l6}�@I�5勊F'�Ȃ�9�.��z�[}�=�Q&��zA�Ov��b���&���#�_u1h&ll�g.��(u�`��,Byto��[�qu5OwS�Õ��u�*mio����'�l��V�����A�ϭ�;4��͇%k�!�w@�gk�1uP!!�M�؀�t((���[��Qꕜ�fo���"�|i�N綛�?���7��v0�G�h�Q�c(f�C@��7Sߵ=0fn,;�8^�̧Ő/7K�˘�CA�d��Bw�|�(n�r

�"Q��(�bH9剕W�:=�L��4��tzQ�YP�]��#�e���t�����Pͯ��碧HΦ)���yւ4�qh�椻F%�Ҿ4I�%�`}� =x�8�-.O��i����$Vc�A��]7
�ö���n���Z�D�";��G3�5W������3Z*1(P�q�x&t�&`����.n��u��jPo�`�`��G�t�/-3��[���NˏO��DaiX++�����4]I֌C�IR��$H��D�ɝ�J��|�d������V�����ƾ�WbK�UVa(��ӿ��Y�?��Y�r�PХ;��(C!�n�r
C�|<O�$I>4��N����&��+� Ö�-�R�gMG���⣕l���ĨIG�þ�(��?`��Lx��j�^d�jKrs{I�?��ut�q�ؐ�( K��gء�"�?��u!K	�OX�v��b��o�[�4 3Š�N4Y)��Q�d��6��t���hh��!�D>�}��v���sgntI�	Z6m|�N��$��WO�������,Y�rs)��BJ[�í%������k%{O�w�����q���Uo�㵫|�j�z�E��Vw��k+Z��{UV<U<�n/BU!�NJ{�T��E�{�0X�@�]Vܤ�?Ni���`[AR	16�>�6r�R�~%GXБ��cs@� L��0!S�_N'h3�8�@xn�2�xL]sYS��N^G�+�.Z���v���3������:�:F�X� +�� /#����z�u�͵�R|��@Y�	C�-�e���h�L@�G���������)C��W��SH�# ��t}{:���3���I�|�ӓDK� ���T�9�Z
-�'���J�7(q�m�e3?��._djkH��t�J>(,bq��R��C�$��^��f�g�/e_�o�����HT��f���<!�dEc����5"$�a&�����I~ v��HS?ܝ�S�����z�ݵ���Qr�JbՍ��6�b�K[6��^^���w�w	]7�ަ�e�5Ʈ��H��V�\���)�6��ܛ��.�)U#��)	X�1ߝ�az�N������]q&.`��r4{�����J�:���] �8M�}_ �c���k:P�Xz�A+��l���w�!%����G�h՚�hB�b�=�)f �6��F��F�_�Ä�IB!���-cMԅ�先S�E��eA�I3�U��`Yy�7 ��u���P\�cq�����џ.�fвҡ��:l�z�/��gӨ�1'�j�RR�{�K����g�9��D��KV���W�vE�ңuh���	^����@<�����w̤�{`�,j��_�pa������)�ā`�)R;�>��A2�fg��X&���z��E@���\VR.=�qE#��&�$�v�U-\c������7�2	���^+��С"otIVY����u5'��ut�f���E����񥡼w�{罞�ʕ��b|��Q�?�:O�
w8�ד�%�����_��C-(Nb��g���{�����w���K�e~`ڙoA���6������|uS#x�������=xor�$YI���\٫��$9�U;6]��c/+HY�G�5�-��Q=y�H\�:�T{���b�^~�gt�O3kk�f��2_9�3��I��#O�l_�5�7��J���]�aѽCb�p��?,2�Ux;��֕=���-L�*q���� ��2/�=j��aP$0�,��<t�#\�3~�j�^�8
�W(�uW��d��r��1�d�K�. �����?��l�I��o�,��� ��b@�l���_pcnGi��6ku
����f��T���y�;��G����?�~��Ӎ1l�>�8#w��ђ�5�V���������������
8�]�*�����5p%�va���~�ω���D�mԦ[C&�h,ssb��r�O��	�"Њs��eѸ�I|(���g~(�)� �_)-n�1�=�y�=�Um�KJ`�!�F-!G����奕��Y
����3��g��l���LERZ@�9�'�{��ܚ����,4��Ѫ,���|Ӥ�d�~�����ђ�F(��D��(��V/�_dq}<d��}GԄ�������5/�-�3G~�q<}~ҍ�g���ߊ������{��ѷ&_� ��
�U
��O6�:��6�d�R2zz����g�
$�nH��Dg�{��SL��3Y+5Cx��2?޺��I�/{�,�*v��5�fJ�8��Խi(jsn@�V�w�45Z�m�SK�mC��͵���l�a,�/ �X�:y��6�-�Z�N�=�}�
�1�?�(���B��y!0	�.4�=sIp�?���������?�k�FMz{T�ۋ6&�9�P�Lj*iuHX�\?���¦��GM��6����a��K�{��]���:���"u� ~f��OړJP��Y<���TB���pl�������
�Q� �/X��N9�
l�Ѿ�[�#�4S?^�^��Xc�(�ZN��V.��;��2���Cu�+�hB����O�Oo �і�Tm.�xN�Jg8���7������>[�@��}w�.��.��L���$@��`w�ར7u��� |���=z0gc�I5�E󠴲�t��c�F�:���dm��`������ .%����lD<�s�Yݤ�������r�,��W�pl;tv��w���Z��Wz.�fy�C�v�zĽ*/�F��Z�H��B��h�J�x/��jq��#�9���ڏi����%��9�I��Ko����Z�ï��a��t���2�{j�h�J�Լ��w�{ �)VE��@�T�OiM=���?�y��a(��!�Az6�J{���� 
&�E���.��`�\�� W��c���fGZѐ��jk�,1��3�T���,��g�Xw`h�@�������Y�n
�/��Ӳ	l_%G�ϖz�7
7����}c�9-5���׍.��/��Q`�b1���Q��z"r���3��f>�Y4�����5�OC��/�^cj�{.&i�a�U�O�g>P@��~.���@V�h�yY����#w��&V����(~�������q������/�K��s0�^a���,�(p�󟭡%�ôJ,��5� ������l�?�v�+~.[��T�wuޟ��p��~��o��{J�9#wovF_fZ��M��zK���W���t0�V(v�o������_�a�UB��|�3�Egȳ�m��I,��Ȝ�b-3�U�m�M��"L��%�4o�M�B1Q�T�
O��@���w��e��4����X,M>b������V�0E�Q���15�@�����吐��ĖZ��%:��ɷ�@t�V��!8F�s��㰋��er�7d��*�i���~l
/aM	Ռ�n�8�V���MbK�&9� pH��t�B��0�%(o6ku�BG�}��L�an�-]�4��4[k8C�	��l���Q�^n6�NZ�P�d��j��95u��l@�{�A��J����iB��'hX��'�%�K.�s��A&H���X���7�b�o�Q���K}�/���YG�V������/����|��S����,�ܻ��/��cyR��� ��q�֑�LsP�b�n�s��U�����ʼ����y9t��NO���kJue�( 'L��F�qW$�C*Rх�y���KW��_c?��:/"ۺk"�9�����9�ǅR��pz	�L~=��:Ŧ�n#�iEg�*���<��G?(�R�m�O��/=>/��M~�{�OCy�E��N��x
W���Qݹ���Y���{�3��3۠�I$N$�k�S])U w!g�[я<
��Շ}�����Sne6���4_�"����T4߃�
w���/	��
Zw����g�}9�t��ƛ�o�{m j�����ʦ@��S����Tq;m�.�ٻ�qy2�߁[�;�%
�?"XN��̵ώ�>�r]�=��>�����b_=s
"��	
��R�3����i������&G;�G�i!uBA��3ʡ��%]QE'�.��n+ʇ��Ȃ �~�!���[%��$��ʷ V!����q\��%��K=��Q�L���s��^�/+�u
�?>�v0;�.�{�+0���Y)�]��צ�T%v�җT�s]� �=\�@yj��iR�%�:��J�7z��a�O2^�h�Sh���;6��Ġ$�ޯ��Y�z`���m�"����Y,���!p`@��Б:Ј�%$�cOk�P�<��� #�Ir�M}�CKX����GM��X(	���Y�.!���֩�M)$2����?�JWs��~^lG��͛�	9��/�9����ĥP�|B,��օn��{���>��\,�A��!pٕQ$66��k7�!��rU�`�z3m���,�qS�9�#(���p�K����.����Ӂ?�c3)��&t D�� �K�N�cm48ƚ_���z�}^�2�J�����HA��(�[�����4��$�dv����H�Rݯ2���T%B�zA��Ԁ�P�F=��c���āYf�d>�i���k��:�/vg��m,��Ϗ}Z�&��5��#��ϸ�2�.�|4Q]n"���; �/�u�����ij��!�&ƣ�D�S��|մ��v�ʧ<�աԙ�B��T���v�AxC���E��U�Je� c�ҍ9����[7�'�F_[M���7�?�l�kc���p�Ѓ�Amx��#SK�oN5�\D��O~���x~�b�I���f�tq(��q�媵y�=F�W�1�{A���lo>.M�XG��fs��rxq�8�n g�GIB�����'Y�4=�B�/[_�����m�7@�[�d���KL������O֛� a�_�|��2@��:�C�����K���l�9�N��w�iM��R��`��K�D��::�3�2�HI�b~� p��.)�T'g�s[�x���fd.�九��z㣰�fL�C��h�>���b����^�Vہ���_��U�=rY�{�Z�v}S��}WjS����ͅ���)"�(i�',�����1#���'F�Y�YiPi4?�j�SK=d?��☱�a.�V��i?�{�r� �A �=D�ꌮȏ�9ZK��M����	�l�>X6��+H��T~�ե�q���K7Ʈ�Y�1/vQX�޿gG�q1� (�$Ɂj9������gf�?����T��@p$+�H� m��X�9y5���ɪN!�
�	(e��hg�D*Vmܠ	�#q�t]�k�A�k=]3���r�s���K�7��5L��їW}������������`�4�=$?'#����{-!lD�������\l.g�022tW��J	[ƃC���o:�e6���H�h�{W�7��Ox0�Һ�+�*dQ���E	F/
݀���.}QSh��׳R��� ��*�����W�{���S{�r^���}��iX��Z������1c�:`l1/�7ƳD�4NO����8iG��`�"�Up��FY���b�(����x��5����"�AC%uw�F�?���f���AB_�O�c$��wօ@92ayM=�f�$[����&a@�ת��{�;�ҟ?:�q`��&6���e�z�$��,�\���'W��"z_�
448���5i]�n~7��Ҵ�B���0�[��ل�{���21a(Y0c�����MۣI烀��Fگ�3�g�D�q-ȑ7k���f��Z�g9u�Xy�%�o�©��=&~�	�2f�7�v؄� ��~��C�S31������ͮ��T����6��{���K�ng=�˨u*}{��y�Ӝ��f�_�EiW:�x���{�{��XlwU�Q����&�.��/��	�����t��"I����R�<bT�����"'�l-�8	����R-9��Qn/٪?gF-�S,]�eT��:4+���W�jG%<���Á~���f}�6��r��H�+��x�es��++�M�_��H��UЉ�.N�?���OZ�fe^����\��Ѻ�7��ͅ�\ř+�xS>�K_���l|����t�d}�����TY���!���[�˭����-`O8o�?�Յ
��Ga�?u�˷;����u{:��`��b�M�������x�'�"?[�{�ÉSA�U4��}�#��Am�X��Q�X_�b&=��H�����2�VD�ܨ"�����{K@<� S�ѱ>�j�=y�Ja��!�t�lXyC�_�* (�@�1Y���示a�}�p�<����g5+H4���{w���}>gGek�����p<�&t�8u�Yb�̒�V��UJy/����E��x��(�M�7�!���%�r��;H�?�%�
�Y`�	N�� ���a.�	~O�*�ʧ�}���&ZS�]� dhЦ��]x�".��;5S��Ţ#�~#�ȿ��ĉ��)�X�X�[=<s��捖i�!:��tά�ʐ�&i�����/lݦ�p���osbZDG�h�H6��k�����r�W�?b�5m����[*}R�"��ֈ���?�<��J�X=��<�:[�w�\��X�Җ!�6,H�*��+-��xjwz�h Ý<��ł�x�����r�FE�Z���XR�rs+�a�Ø&�\'�JF6��L>���t�¯�(�x7є�S.!aS�pyT�"��[piWw��l�/NTb��#y�9ʢ)�T��)�(�X�����h���^�p�}�7r�S�3�2�^�C���_x��g��a}W�ͥ�ɒJςG��4�%�Oa�k	�Vdr<�8-կW���5��!GoXut��S& fS���!5qlr�=�"/����5����P��D�PxL�)~}�e�~z�ؠ]�'��SeC�XՃ�,TE��ӝ���Y䦢�D��qZ�J��i-��@:��#����Թ�X*�|)�?�#�����8%���	�G�2A6�|�򯦁6�CIr0����ƕʧ��5 �Dƃ�_*Pk{��x#��E�#S綕o������}��I�&���=	�!!�}���2�c�K.�mDZ��ܒT;C�Qi>
���?��pq�ç}�%����cY^:�A���WHD#�C?�l^dn�0��?��h4=Q��-ۣ#TT�����,�R>�3�Z*@6��b/<(����0�N�\Z>��=�Ak���!`��}QDB���A6�2� �$�V�b�H>��T�oɪ�O�a��-��)޴��W$R8ׂ� �o��L�<�ʡhQk������_�%$�<��,�u�ߵ`�  8:&6����%���R�����N�s�F)��F�o��Ec�����{|'3����g���"���M��P�ET+2���U���씱��#���`�ԺD��/�ҝ���$�Ph�ėmj�u���z������QHS�J�Ҟ)�L��� �����l�KP���ι��M����;��&����Y��-tpAY�(y\WI���#R�5�s����*���O~��fc���U�Y8�����%�l_=�`)�r�6�OR��3��������& �?S�V��IZ��.�-ʨ���|xi0��=z��(�X)o�ڝ�/5(��%]�r�W}������$�����{ϙ�׮��i��"��"�
���v<�')��y���,�|XP�t��}E��xwO�w�pj-�2;�5x��=������9ъ��Z7Q�����ïq�rUul�	�N��A�UxOF�O��������l��Xc��m=�9ţ��޺D���!~Z��m�E|�)���YX)�����u�r(O0�Av�Ks�Ĥ!\����/+/?���p�u�2��Md��z�
y 1?��B�kS�N3�>Mkj�B�6��'G^WJ�����?�o\<=�XGX� e�6����6�����5Vwal� �İ��5��&���cuSȹ!�YB���`#���zu�����,?y}�l�;Oh�)S���tr\�x^�V�0n2l�q��f�e"���W��FQ������fߓ�A�8�~��d�o���9��c�#b��QL�/�F�j�#��f��I#���R�*j;�#��
���8o�4��������@H5;��߻�&j	��|q���Z��7'.*_��'���F8�=s��}���W,�l����g' �|��+71�dîY$�� ����Fr�@��ZM�;�@aq�AP�K�և_CK�m&8+��_u�2 ��]��c���󹘫-�Q��AWͿAa��$p��֝��n���p4f��=�z��"/إ��n|�iWɿo�z_������!�@N&fvM%�h���ӝ�w�����߶����'�"V�'�ޓم��N��6�^������qu ��f����c�fr~�R�`� �_��J>׮��q�?�gy�FdB7(�O6������Rb�C��P�بf�-�!�����W�7-]ȿyev^�=R�O���r�"MǇ\Z����L	�{y�]r�*�d�[��w���BPH��vx��H�I0������T��u�\;�M;SJ#��B�A��'V�^վS�4�t/�Hm��mw����߁���&�z�����8���j��ZN�����(C�NZޫ�b#F�q;�ka��+/̴���.���)Q�_�� ���%aYs�du�ϓ��+/m}�����S�����C݂ٶ�B�Kt#s� 1mDU%ۧ����ɭ�W�Q	s����Ǖ�k�#`���h�Oo����O
�Jv�'�*f�:���6��9��~��pp��T���)��
�j Tn�J���q�SǔD�r:{�n6��m��Ed���o��0EF�#�&�O[�����[W�0�0�6�C���@�u��*H��nl��o(̌����d���SR�ϵX���Ŋ�".��U�aw����X�ב��/��1h�����G4�"�/�6�8��xO���XO4���^��FC��4ȉju-UP͜@u�o�=)��h�S��9m�P3,�NQ��Ėޢx�c��#H����n�=��fZ�{Y�^Xiۃ\���

"(���C�Q.�
3�o k�W�mk!tO���?�Ghi���� H��o���9��JKQǨ���2�l��J�}>���n&t:
	�Z�I�o�|}�����K�Kc���:v��zSY[�d\�f�MK@mP�Rt5��(�8�l0?�
d�����Lx'�$�M3F�T���ߩ\j�uB�������=>iQ��L��mg��Y�h;�#�,ӥi��(]�b/l��o6��%	�7N+ P��؃��o��J쉑�}>�8�/4������Vzޗ�ϲ�t�
=�l\���c�j5��k���v�g#��V�	�7�WГ��6�⾿�{~/�	!�WW�$�YJ�h4�妧�#m�8Π�����}�`xvp}IR��P�?>o�M���]��kk�;������������A��5 ��T	��(8��͕6����a1C�lx^5���{�6?f�N�Q0��ķ�bE�'�D"b����)n�J��WO@f��e=I|BZ*�����XLLHed��b_'���P#�n�dA/_*��������t�N�`n�Ю��PD ҧA|I:�	\��g#�H�n�{~�Gv����������V*�ֿdk:<�jA\b��'�%�PU�P[�"�D>X?R[�u)j�=�Ld����������Ud���k#��[��ar�2�܅�LSBE�5E�<��t�%\��#D�~8���C1;��S�ip̴������6��
ެ3UdZ3�␒��5���6V��}E��>�⁎�#k\��LS�#��R}�Or3�9�p�.���-����`ӳ�����Ed�z4��>w� ��r��,��b]Խщ�m�?	q��D\ʦ�;��E/�po(c5܌�#�ʥ����=���l|��eF1*h�v�A��h-�C�z�I�6��al��9p�x#��W�{���lf
�D���}<t�y0�/����*u<Rz�G����N���n���%<	J��?RSL����	����5�b1�C�K�[���y��6'��)�(?T�����΍�Һ+U�����iѷ.��/A��R&��\ՇSƳU��NJ����ĭ�Z-��w��(z y�'�LI6����M��Ň;�Q�&ɨ��_�Gׁ'��?YΒ����{��v�7����.~&�IT$� bZ�ҏ��A�Y�b��r�$��̬
%_�ܤ�QǑ��(�Z��m-�6�o����X�o��H>�|�%��A�oE��g��RYZj��Jq=ɔ겂C�55q�	g)�w����G�0o��eQ$Y�ƈP��&�6v-d@��j&��X��/�o r
C����ӌ����<�/L+n�*+[x-��t	.�&�f)���x�̰�����S֠e��= 5�͕s������98x`�$Yq��;0	�ڍ�),��t> �D{QE��l�8�zn��9����{�W��*�T�d����p�]U̟�����H�� 1q^B��R�z���c��^g��!&Z���f ���7av�:�_)�)�<�L����J��L����%t-��4�����kR��H�̋�b�N(���o(�,����vAʓ�]�pk��8����o��������%E���ǮOx'�R����)VXM�|S�����L��ח��ژ�>t�㳠�E�ͩl	O�v:�>�i�K��f���H��pmm��k=��A�E���?�Q��Ϳ3�k�e!���5�zSc''u{���%S��D��^'�[�CˢK|�n+��A畓��ʞ*	{e�1	���5G����|
��x���:G0���)�Ϣ*MW��y�d�9A[R+�2��W0\��U�����Dg�=RsQ�z��63󀔦k�۸��g7�1R�_�9���C���I���H��qw
|NEf�As89������.C;��n��Ǿ{N(av��*��F
]�)M���s�bվSgD�!6�� �(��n�dK��C�p���Q�R��;R.b�#�W�R�j�o��I(���'�C���	�7c�sBc\Y�1��5>;x�("��}-"�K�&��e�R �t-��S�?����@��ϟ+���~&NR�]P$h�F�f���T1�W[�f�X�����Hv{>��$Ob�� E1#ԣ�@9�;��O_�&j�Y��E�jK�C�#�7a����Vd� �m�'�Jk�]��ᅫ�؜���?��F�t9��3�·X���_�m�� y)M};�d����\Y��X���a׳M��'��b2��<A-��ͣ�ކ�j2-�?����������"����خ���ȇ���ݟ�-{��$�����}Y�r�C	}��\#:%��|y����fTI�Zl" �d�5>Qol�e��WM�̪t���yV���Vs,C�m,�}K��c#��%U�c��}��� ��ZG���Rx��7��m�_�|�O@�́<K��'?�3Qu1Π�BT!(��.�����ln�hdBa&��<��J+��%ae|�Ϝ�C7�	�:?g�Z!���O�u�@0�s��"�Mޓ�_`�B����
�.F��`ړ��{}Q�9��>����MO�clʟ�{J�-�^�P������m,O.����fv�]i�R��K��i+"����@Yoi�x/�Q.sr��+��ܚ��)�*�V�g�{;��"�Z�t=$R��KJ�d"��[�H�y�����<�1c/�&�Fw����tJ)KផU��6�h����М}:.�ml�guܛ��r�N��ʓ��������VΦgW�t�r춥Tyj*]�T� 0��CS )�r���Ϟ�2|jP��(Z������X���m;�9���q3g�c�����Q�B.ډ�YP�h�ڷҋIƜ��7�������3����oa���q����!#�4��wi�v;�JI(E��օ8s,�<�_:�rQQ�b����1��KV��ĒIDx���@I�����?��pe�%f<o���׈UƯ�;�-I~������'5w�����y�=�,�#�����X�E|���%ܫ"jy��S%���r3\V���y��'\��4�D�E��d�%o���g�i��cTzp)q�}3i�0��F�0�ĥ��d�~ �������gS��iHf���'ݷY�Xe��t�6�����wZf�4���^��ޡέN����� $�[��2��;�X8j��o�zל8�����4��*O5W-_�Rͷ�ʧ@�Pᤪb�fQ��w�q����C�A�iY����9�����Y�ņD=)D?h;�Ra��_��b8C�����|��N�������(WĲ��=��N��V��dUÉʄst�:��m����H.���'�VL��fck��E3�0��G��¿���=`�<.I��P���BJ='������>Q<b�d��~g�������WRp����4�Uw�=�qk��2��p�ø�1�▋IB��7���ܷ����jk�Nڃ~uH�{ӻ�'��ǯE�Z�l.�L�z{_4�m]��,��W@v��	�k3�k��"��/|:EaE�/�y�~a�;�-?[kt{Z����P�q����4~�/'j>]쌿W<H����n�'I��H�s��~�H�'',5"1Sm��2���4S�:*�F�yFҫ6��Q�P��N�/�PLg�%"K/���*�aK39~^))
Aq�\�P�z~��� ��Ke���cH�ս��1,�W����ރ������*�fg��l��{��f��7���q-tc���Z�'�I�v���+�t�5
d�<'��*��H�:��3�g�*�G�|Q������K3rq!	��7��Z����g+�����?������?�^����x�"�%��b:�lHW4�&�4������\��4�/fsju�_+z"����s0=G�Ug���ע
��时��ڌ��;��ǅ����FWe���S��?�~l�r�G�)��9��{����{?��~�!��a���Vs�=2i�N�h(+�<��n�qQ3����Uݒ�an%q�&��G׉G�S����"R$ેd�э�ZU�]��1���w�2�ktOu�7�<�����tb9)
��$���W���w�/7�ňpj��S�]��2+2P��Rp�PS�U��%m�%zZMI�AL���ӓ*��h��^Ҷ��.z0���ENs{ڲN{���<��#���pi�.ӌ7@^ ��O�Ɩm��LI'�����Q���kĦ�]J���b;��wR2�V\!��%���u�x�"���ڳQ�iQS�Ϝ�0��3���7���UU���e[�(�^E���s��������}�9�8�H��C��V������3ޕ��Buef��UW�W\!�����_,[�UK�Z�r|)]�FmY��[+�y�9!�|XXj�*������:WLjsc�as�Clk���=sIqy�@�BC��&�\}��/�=���V:���������%�	pf����O�id����=>ڎ�P���X^�6�؋��6��z��y��/~��Q��y�
���B� W
~j(��M������ʕ�5�����-w)�w��/�gӚ��}'�AJX�d��YJ��p<^p�UOV�z��=�y0ASC8�'<q�Vs�iv�G�����b��� ��̺�MT��W�D���!��Q���[qޗ�u#h�����B��F�9���nV.֩:O�Ec{��v҇±�y�q�����_���ߺ;{6y;�.�w#ɢ��;U�(3�/����_�b��0پJf�Zd׿H�QQ�	d���υ��wy������~y���znu��:F�¶Ս�>�����-�z���/���2�Q��)��:���_�n6R��Њm��wk��|?{ 3y�ED���q3؛�����T��9�"j��ˑ K	��C��9�=酹*z�3~�~_>j��w#�< g��\�IGl��H�h1�bmy�{�q����!&������ũd��$�NX��0��,,C�a���X=-�����Y��$8�-��Q�cp썠����/���}�
��Y�X�6������Y=�:�_r(!�j��A�HNy���<����-Yz��� �2v��~��C@	+3�
}ǫ9��>�bu}��$Z�:��!x���S��2%�4��r� U��H�Ik7�os��ԣ%i��-On�W���5�T}��8���'��V.�UmWUx.18��=��nVS�
�Y,�'���V���4� &Z|C[=7}vol��&���?G+1Q��G����n����B�T��An4����|����М�ԧ�/%i��z�^z�:l%���O�g1#n����<Kݰ��7 �ow�ө���=��	�7�Q0u\�N�V��o0��g\&*�\`�l�j��BI��-�ob�G���C��7���Z��0wV_m0��/R(P<P�8-N��Zܝ�ŋ������!H)�����{�}��9�s1k����f�yFEF\O>���P�@��~3X��k$j��w��7��������W#}��m�����	�z��?=WGP�1�:ޛ�K$��G��k��[�	c���$�8̄��v2ۖ[��
.O�T�Q�N��1k�G=F>on���_lDx��g�c�������(lN�y���O��٩��<7G�-����A���Y�<�R��5-Vi���)���J�]L+л�%����� ���6$��y2��g�q�/ nܝ��4����'9��f
b�gb����#钧WS)��4�.i��)�t���Z��Yӻ�]�p�$=%]��_��>���7; �3��b0��R��b�E*A���S��k�HW��LU������~�p�bf�W޿ Ҫ|�!�٩�a�/ <���滹�8�C�XQE)Q$w=c}�S��?u�T�k�,:O��KY�k5���0��R}`����𹞡W��E2+&�qOu�]�%�rh��).�!!���6�w�iu>٫`��0��І(`S�lY��nv���b���c�KL;%/��3[�-��U����Hb�ќ��T�OtǪ��b�0��W�
p�U��"����.i�}g7B�g��U���˛������.��1�`��L�g�lt\�I$��Βka�Ҷ�gOT\X̴��g&�f9%�ՙV����x��p��F+/�/�6����r��K�O�x�+��T�Ɏ5ү��;u'֐:��+�(����n)࿯\ʷ��^q���V��E�q���8uuS��*{�ϣ��լɇ|�aP�:�H�P�-JJXC��+�N��=3�z��X���h"�|"5�kE��@�����ơ�~�/ P��w�$��NL�F��3�f/C��k��=�O�j,u��?�Q.��Ym-k����m��M���@fw�ʖ�>�uw 2$|�QI���ZQ{��Dm�ݤ��*����A�3��N��3����S6O���-�����7Ǌ�0%O���3�?ۋY��=DXm��l�~��
2�߬4O�<�>"�te��/P�:���='�&V?c}.�˝3��>�XR�A�6Yx��w2�rP�tL�s9��ʶ�(�2�k����f޻��)�X;��q
�&���.���������ߝ焠)�����tĿ�	B'����	q�󾣚_ ��Q�';�0�h�戼G���'}Rە�)�J"��;��d���MM�0�Z�7 W.A���̧�(q$ ���}���ml���q��qJ�Ӹ��y�$�J���iq�5׷ �oC�����kџR�(�W��+�S?�W�5�P"w�N��y�޷N:-���!�,�3P!ӫYS-D@v*_������M�������0��w^��	߬-��W;���R�Y*�
v q����0/0G�y>	+u���ov��f,�9�MH�5ps_Y�I�\�;Ε���c�}*TGܕ��S)��PSh�~���vx��"��آ���lb�PϪ(���Ա�ĳ!�4I�k�x��w�U3�OS/��\MZ^ά�!�Y2����g����t�z��jpZ����6h�@h]�LtT��0(*�c��|^��{���ح���
���G/���W-��N�C�RX]R�+�͢WQ��,
_&i	PW��_��	y'��6�T�a�?]"�p7B����~���/ 4�f������n{��}M:��	_��d���ۓ����G�Gg�v)s�]o��o�iiU^ H�"xha`/j�=��[v��?���t��7?�dU�I�ZY9-�ƌ:�Ӝԫ%������l�� ���.��'л��jO
3�����������Fަ���$��A��2��e�ao��k@MUp��i��
H��^ϖW��;�}�QX���8G�=�(�~Fm

bF^.����L�yM*��:��z�g��@ �!��K�2��g�mՠr1�M�����]l�\1�f��@��?�LW.3�Am�X�?\�Pw��9ٙ��'�*LQ[�s�c��	�DS�y��n�F���*�6��~�s>��C�tx��n�n���� ���P�U��1q���eYP� U������1���އ@��1z���a�ɟ))iG�����E@:��X�2��#k��'�{j��I��/�T6������v�1�<�Ռ��V��S�ɕNF_*^��{��q��_�M_F������h]U
W��
�Ri�h�01pm[v�ir�3Kґx����s�-ev�~� �E���l6��s���^�T�ȫ�H�̨����Td���q���?����)�����=j���sSť�=��;�n�wT޳5:�;"WF<�8gyzh�57��߰X��/��'�@�|OL�CK_�<Y(�x�n�=�X�ҏ��q��Ao*�u�����`�#�7o��܉>�+s�e�v� �����Z	�	$HεN8~�QurFEV�a^ٟc���?>� �A�]�jvRT)��ˉ�f��3�pM���Ê.Zȇ�y>�_���ІՈZkg!ڴ�%헏^,�/���A�O�H%�l�Uz=bd���q}�'Y�-;����ʗ�²��VSX+]k�����_Y=N$�f���5[U(Nh�| um[cҐ��#�	a�b��w)c�q����e��ϸu��}<ڙN��@�G ��	s���8�� �V,L"?��}���U��~�8�h'�$��YyE�i���Q��^�g�]�Q���[�H��x�d��$
�U�o(����"�|С�D�I����Y�X��4��c�{�ӯ��������~�	O�=ۚU%�V��<��y'���]HVDN�y ]0�!�$fEB�2^pC��}�|f���WT6�R��Ņ� ���I$�J�����K�OY,ȁ�����c�V\�R Ȳ���m�M��\���P5)��i�&|�������f]��&�	��8cJ�'RK5͂��:ʟXT&l ^C��K:���)g�-x�C��䞞�Å�R�X5gN�`����4��5�2sfu�-����0���4>?z� ���i�|�l1^ D�߹�EV?��D3�DQk���-���,��+�I�N���E�_!j�=]/���1ҳ�>Ϳ���EOr`���]\�\{y�<��(5�'��on���^R޽���yT�ڝ���(@e"�ڲ��JR�[���>$��I���9�v�')N����{f����/�ԍ��й�S��ޒ��Im�~$:*!�
�9B)mc��\��i��f	.B���T����YI��X6�QX*n9�b�إO�>w��Z����I������7=�0��\� ŷۜ��v��7�B��$`�bWhvǽݱ9���.�Y��e��J�!������ ��C�J�n]�넕%Y�#��@�kb�1�I[�����Wh�$���Ę�@#VP��z�e2j��5h�Q �:�E4i} ���k��Ϧ��zJ-i�K}��y�7�\֡�L}N�nM�U&�����)5��þ�c��i4O��cy.��D(��7�|��j?1�[[�}��o.�H�^Zm�ȕ#>&��g�o,�<�3E�&u���K�K�gfQۨ9���":Mޫ�,x8�H�<��Ej�B?�L�@{V�2��2t0�D^Ԇ�Z��z���n����lmR:��]�ߖ>��Cs8���%�w�5��H�1�M���Bg8Z�����&?����T+����|�];�`�8Ayf=�|D|}�o�x��L�+S��|�L+���r_�h�e�q�{X��ҁk�g�2d?|fg�{�6u5��~.I"b1�buI
�9ʥX̓�u�	?1�A�/�����	@�I�hE]C�eaA����8���Dt���Oe�U���jx��P��z�T#�_�kJ'y�b�$<$'�!DV,p�aX��s �����Z��heJ�h�ɤ$6�i�S�yB��8<�6��ND(ʈղ}yR٧G��C���gp~U�E�/D(�kw�"K���AHZ>F��Uۋx������G�������� �����&Xg=��HqBvVkP����^���0N+�T*Y���O�[��.�ɜ�eq��2�RU�c�)~�1+X/�q��*!hWm�7��H��-o�$��ʮ�`!`K�O�K �y��T>JbE�[��:������[	�����x�E�ɮ���)�~r�B�����مO��W}�g2��BkK]�:F�eY*���/�����Svk�f��)�֥���.���\W�KD�	}������t�^��o�eݣNj(*��`:>���N���Ѭ��4\_��ք�Dq!Fv�u�ܡ�J�MTy0�/�v�u�0'hb��:�M0�2�P�	{5
������mq�k�_���!�G�p��/-M_<`&�W��ç��/G�0bڣn_U�1.bz�ӽ�,#����YJNJH/����+�ۨ�{c厵�2:N�Z�͸ˁ�n�1���d�A�T��?�Z[A�&���������igk��m	|�jA��y�{��X/O��M��qɌc�Q�@�`L�"s��F�����q�1�v�Bȡ:٦;ܦk�2A��<2��\l&��y�wնS�[Xk�t��;�-Uux��q���֒�bZ\cc[���b��:�13�T���Q��DCX[�O���*q�Tv:��xR&����p�sC�X|5���Nd˦Ƅ �q5�y�^!�z��
LAriTƻ����Wt����}n�����4�f���E�Q>�Z�7Zw�������l�΁�!��ԓ�YM�=��׌o�;$x+* $�Ł��0m�o��s��T_���I���1�����7�IBYj��')��k�����K��7e�]|�����q�,�2t��G�q�G���n׹FQ���m���n���[�ɥ�ef��|�x�1�>_�Hwpd����ޒ; �;���0�*{���W�@*eG0Ҽ�V/_�3~����ӛ$��.W'<�����^&e��y
.+�<�^h��d+jˣ�Jη���Q������ѮQ�*\�������O@�|���E�7��?���)��svRX=;�xIE�G�� �]6i%��7Q�4`�P$�����?�GO����G��~/Td�Q�fߎcv�P��y䆒�\F�Kh�������84S��Ux�1��7�z�)'������j�(V'�Mɻ�ep�E�~���.B)��q�Kf7ظT2H�H��><�|b�M��_;�-e�bC- ��д��xT��OM���
3�(p��'�T�B��bySm��G�.b{��̎�Ic���f�%J���{�W1�P��43�>� �WI
ӆ5Y󩈠'�	�Q=|���r4*ʜ�fI5�E�oM]sD��r's��G���n��+�X��.��S'0��CRN�Ԏ>>�Y�y<h�_)E6:/�@��E�K�qN��Q��mи�m�d��Wf.�t�z�8��g���4ۘ������mTUƧh�$u��t������=����Ŧ		s��H������KN����89�R�P�==�_pʪTf�E�d��,5��3z�Z�--�r|s���.b�.N�$�z��NM<ǒ�Yk�j�?�M=�����NL���Xe�ή��ޞ�[�k�7��]����_y~?��^s��r�(�B���D�( 6D�M�a� 9}����4���U�?��u����L�&	�YL�(� �ɻ
��/֔�YD��!�<��ˍ#�]>���
���x��kآ��jv	U�7��rk�<��.(���8k<-t�]��,�"��ʉ�Rb���p!���4�H=pr,�goo�)Bn{b������)������~���t��j3��~8�|T�V��F�[5
�t�y�N�#��m�my�H䀝|�e��k���Ğ4_;B�mi��g�u�;�"�eEx/�F�OlbkKEx���ޢ{e&1;��WPq~���;��F�3'��r�T�<�̴Wq}^PGoO���Ȋ�1}2��
!.�:g4 yK���,,@�K�ZZ<�@`�9�X�3���w��a`AL\yy�f%�y1�:P��ާ�!
���8W�OR#�(S-�:;V����O,AF!�\���� u��
7�&o�c8��)����^�V�4��  �#�+f^T��k�<G}�i�[�I�o���i�������u7������ZĲ��#`E��w�$#!E�V�+2O�d}��&��� E�ұ�n���J	S�eA�}�����\zr�=I����6J;���Z3�����)z{��A����'�V�M@(T�W ��������Q%,�X�V1��i��MJ�W�dv`�2?ؾޜ��*}:��	э%��Y��֘��A_����c�܎�܊~��͇�L�^"�rm�C7�6V��X/�L���Z��f�[e�!���bfF��C�{l�]p�"=���$ŝ@�:��C\�����~��;O;Q\s�6�h,/V��Gj�cпPt�����9M�ǅ�x�s=�.�M���)��%����#R��Z�=���]*��6��@ϛx6�k}`&����T�+Ƈ��U,���U�^8e���s�Q�p�t	|��pes��9�$eu���}���~Tj�?�lh�}�8T?+^�%"� ����o�[}��u�^�b�p��TÄ�Ww&�/)p/�a�#���鯿�'��x�~![�(Ki.|�PF�:���=���h�w�el]{�ջ̼M;���2�d������'��kJ�,v�v*��f5�b8ރ2��<�n�8k��ݴȌb�������5_� �D��=*�����,�|5��晦��~[���#b(���7�&�wf�5t�S4;:�&uYz����#��ɍ*�m_�+u�@�DC���S�����5��+8Y@�۽3A���hd��%D�k�j�h�R� �7�ο��t��M>L��xm���1�3�̝Q�0r5M��34+�F�,�g13�u3-[1���2�E��z��ukp����p~=�kE�o�E�ƚ-�`��H`Aj2�N�R�/�9��T?���n� z��x�U�}v`��1������N<���;K(m)1�pl�i��<�5��U�.�=�������F~�x���}����\^V���X�w�t����yc��؄Î~�o�F�k���q�V�(0{�ixO�(5����7%��<��վ}J�?i�H3$Ghn�jf����9\ �w&9u�P/��c{����	8�
3jEC��t��G��Z
lG[5�hŮ�-���=��4}~��w5.�G�6��S�~�]-��~�&F,��$�I�x@�=d��l���&;��#k3�~���T5h<�x<�R���>�j��,�z�UN�)�/З"^�	��&DX&�$�T�Jh�묈��FP9�"��P8�l/������}?6�̍��UQ�kdb�����('�DK���վL81�ϛ`�3�]2�}~��O�pl)������X��4k���^צ�-�){+�9���I+�^��9-�Z=�#($b��D`��$X!A��S͝�6��:z'��u<�.74�"�F��2S(�w1,�@(@F5���ܵ�`��@S��OT���Mվ�ĵq��ڨ�W;��мOc��@��L��ց�<el��I��+�(������D(N�~a��3����i�'�;�fo�;�m�k.:����I�<G��p�L'`B�ն�:j�!2x�-��ǜP��%}��hC��έg4�VُC�b��0��"�΁f_�	���8��Y������#꟡��م�)�M�t�I�o�R�B�'O�6�yߙ�[C9�> ^1��	�N���X�{�sc^�JY߸��.d��=Be���0�p� �+I��(V`>����k�����6�u�g��\ks�q&;�>t�G��À��l|.s�>#��	Y$[�fE�5}m�4�[վ*3.�Iyx���9_��t����t��Q~�s�������QQ�<�����(w���1~�n���C�䶃������َǾ�\�Em��dFU���p��8�Z�
�1��X����,�"n�׋��/פ�[r���A@E	�lv����z\m���)�0�ny�Ӻ�
 a׺#�"��|��8~L�"��F^<�@��I�Q��~7u'n�_(��z}5H&@�V��A��Klpޚ��V,�.���)���\L~%��H$O6�f]$���ٍv��V~�_�f59�b"W#���ƚ�&��P"jྊ�kfA�c���2�>;���1W~�&E<�35z���aU��ꖜɑ
�I�-���²;�;����jhi 8s~�[e�9���(��x��>�W��u� -h'1���Y/�@�L3*���q�Agy�k$F�{���랣�`����*�f�������_�W�f�o�AZ��Ȫ��,ۆ_G��Zꭏg4	��/��n	�Q�Q� M��!�v�D!�x��X�o����f���#F�
����b��:�D)i�`���^�9�_P��;Iv!�|�6�a�4��y��_5�O�3�셿���݃sMeΈ��I$�t�Ծ*i��)����ʻ~�U���h{��dq���M}di�N'@_9'Mq� TF�x�`+�x5�ڹS�#�o
��,���y��_k�2�>Q��OFa� ���.��9�2P��4��h�3#jDK�?[+�^�O���ᢞu����S��c��������cv�@�=P��w@5�-��s�h��"�����V��ͤq4w���g�.~�iZ�%�����OAH/�c���|w�CMZ��4�Wc��� hY�(��ǖ7��@��Z� ���S($g1�bt&�yd�S��4����ّ>��������`��dp�M��oL�X9-+fM���f�7�#���?�?�wd<s�h[<H���>� ��\��;�����Z���W�����O{��P���A࢞A]3f�֛���o���M��#�*�\HΥrķ@gS���FY��(�_f �'�|������X5k{��;�CL���A�Gӭ���0�D���r Ki*�_� ���yx��h<p�G �6U{��:%J�&���	�6���^�.%�?��G��!�X�������z}K`pvV �0�[/�a��+7�x?f��̵���Er�.Z	'���?��-�5�Z��=r�����/�#���6�Zt7T�[�{f��5��}�2\�оF�g�vyn,�r��ڿ�����b�����ē>a�J�7��[#a���s�_�Ü�<Y����k?�:luLR�虏��8(�u�&ŬL�?�x�(�9Ļ��2N���DX�D^��6F��0v�H/Z�Sl�`b.?:�UZX�N$�������>`�C����kdh�S�2��vQy�2�FW#wb_ x��fʌ>WW[���F�-�s<_�(?1yW���N(Gnь�k~�rw��vհW�2\ Ş�4v���%V�s�88�4}�~��~{���#XI[?�>цl�����C�N:d��՚��	<f�eV����g�����:Y�A&�Y|
�ּ��M�YQ�9��^����q� ����'��Jvq��H�e���զvRq;z��.{��^x�%'��,ƍ'S����e��!Vt� �ڬ���%�'�R��x9���U `�&�����r�R!e8�=�$/��\��{;&��#��\�/�f^&���[D�q�g��
?ȍE���G��W��[�D�n�s�V#��U��P��I�ͱ���V^����LQl�=��"��RSZ�[���84%P+��Ǔt`�+������$��3�B�Ϙ��`<�'�g��.�@�����!�Z��gͪ�f��+�������;��r�H�Z�&��M#���{�XD� NC���B��b��AT�Ɲ��Q:;j�sQ��,�7�_��
�J��R��af��Y��e��G�RK�y�e���BV�G����4�RaP����2�ҫ'o�.k�ñ�`�S�����Ӹ�Wr�3AW��D�YL|O���f��0"{]�E��3�3|�u%��q&���	��<���������^4�{3�۾�)��#��	�)��3ʇO���d}�6�~X�A�D��̌<w���u3ᥘ��F�(�&��k8!��j�B
�{[�'3Emn��6����Z�`���ٴ�2�8�<�-�oE���q+��6����\�|4�S�Ԥ��JFTYl�2� xٿͧG�9�#pU�$��ě+��8�&��JTK��~l��ԩ��.P�2F�ʭ��W��d���h|߰s����WQ�&VK ll��y�CcY3ܐR�C�H*��F��<^Ҿ�x��U��_���d�=��t��ݶɶL����@u��*S}�k,�?qϧ�f�ݿk�]�n�_E�����-����;J{�OT{o�,����+��l,�z��?G���F�/�˹<���mť�61�;_�4���J��ĥme.��Ե�ރ1��b*S��F	O��o�z>qW���Ű�/����=�_�f�������)MA����k������)}�*��"J,R��&e���H�J�z�᧌��*��;�!�%Kg{�_��,;_�.�/�#���s>��'���BB������T{�q�j�	kl�5s\�w��d�J�\��0Gz:�\�j��6��]?)oi�GJ�n#Kt(��|z��;h&�-+�i ���@�<,�*�+���D��>Q���l���Z�]��-��j_��L���X��K��
�i�gn�Sr�5�Y�hdሚ�5�ݒ�jHz���G�vw�>��CO�m����:1!PQJ~h�,�f�G��'�8{v���\��s�`�<y�qCfUTyn�R��;��f7�rEj�߯
9��6�n6��u��b[�m���'�P���#��X5�1�f�f/��X~�	�
l��~Ym����Q}��j���=���&�#d���o٬C��=֌\)2�������F�󬘄��%/ 򅵼1K�%��^>O_�l#��S��ԯs������	k��z����ײ%t��')� P{>�9#+�� Ʉ�k�y�n��l��q!U^�[�	��CN��-έ�CL���)�7xiT=N��~d�/  �m-4�ʭ���J������T<�ʍW���;ݔ�\�ʍG~��1��T�d���i]A?����2#�߸$��3�x�Q+�;���lםqI���n\p���󱶛���! �����$��ġJf�v�*v��jw��堺
,RN+���{�\�qsz6�9>
SN<s�z��~��s��L��r0��W�0�� �D6F������x���:�@XՊ��������(o-9,�~��K2.^�U�D��_Q��>�����)����� ��K�Tvg=�ld�Z��W9`5�.Ļ^|d�<�z��7�b*)�H��3�T!�����(��1�!?�Z�����/*F}ws5Gr�/G���a����R�t�����s�of�J��U'��w�u�u��x���R���� f�N�62Nhc�#V_GA?܏�a��{G���M�L,��"o�٨�۩��-世�x&�_��/|U�BZ�	�%$�^ VK�������7�d�3�Q�Y�t�vz�!�0��[�\�`����1ԫ�ͭ,�p�!ǻ�j��k��oTZ�����0�B|���S%�6�LC/ 4�����r���݅XK��#�H�=�yv밅Q���D�,��"o7�F��W�^��;��Νy.V��ͼ=�	G\�Y�����ץX���G-��V91R8���{��l�ra�"�w��(��f��N[����jSy�l�BQ�t#�P2ݮ> ��'��:���K#������C�➶�q>�a#~;��#�k�UH�Z�[RF�����/��x]|����6v�4_ Dj�6p6%R�\�����������i�>�xy�:E"��w2�Y��T_ \��5�{���f���]����2ȋ�����n��,"�5��Z�����d� �aye:qܘ�.w[=�Z�=�:fi��s��q9�P�ӱή�brc(D)���H�)[V1���ʳ���ԏ�K�t��O����������PU�WJ�vk��`Wb̢-���c~\�f(GP���R2hW;N{^6	z7���� �g�ucw�y���I������T���f2�J\���g��� f��_$�wIߕ�%�s����@��~������a�,,6(���9tʕ�$@�>s��xk�cXB��O��KЫ�V?u�����N��/��?-�֚>_�>���7��F�3���Fj��Y
}l�>r2�8=�q}O��	-l¿����Z�.���quV`h6���$p��J}��@����0�|;u���¥�~�������c��|i��O^���(g.Б����/*6x� u��t�jg�(E��4�1,����2�\c�]iճ�*5P�*�ή�`�cy"-��#���������9�@IY����^��/�.�wKn����Bo�ҫ�.6U�e*�ڔ�HX��[k�Y��7IS��
��'_ ���҈�K�^]l�����Ei�a۝սY)	���27�Ɓ�7���!��c���b��]]-�������"jE�M�a�ZtqF?�/Juͧ���Cg���u�0B���?�?��\������<oɱ�с"܏�@���RT�K��%�����ڒܑs��� ��C�Kh���rr�FT۾�K�*dne������'�c� �7[i}~�v�}���{�Gr�+ ��'�Q�3�V_��ѳ+y=�р��i��6��2���0��D�v��,�e8��,`F�T?�=u0�
�1۷Lkw!��h��dy~��D�(Gz��<Ŕ��.�x��M���f�u��rF��]5-*W�.��	���� ���;2����o��W���NR�m���J�uXI�J��]�&�ݟK$QmΙ�qG�{�so�Q���4
CSɘm�ER����$i�rT���_����.�g�R8UY/b�AC�y��z9����L��������L K�
j�Vjbu��F[�!�V��:���/��D`"{ �c��~���4�d�K�=�`���F���%yh�
�ä4bg��Q�Hg�M8���Ff3!suɞ�LO��!�����|tղR\J/�q����B=����4��c#�������]m�Vv*,Ѳ�eC#���v7qAXYMTs�Մ1Ģ�>���h�r����&�O4v.}������j�-�])XޚnJM��`�e;zU��4�����+(��>����}���˨j5���M+���r>�2.R��+�@�r�|=TG��8~3��٠�LE���ß��r(��֦ŭ�E��b���??Ux�������QhG�9�!��M�	��H������<�[$M�#y�4�����y�}�3����-9�'�噳5|��߬T�[F�s̕�T��:���ƒu���?&�}��\���:<F��8��d��8祙����[��@JR�&�ڻ��@R�2� y���.�q��V�v��TeR3k]��p�q���.�-Mq9�d�.7֮�7�j�A/>A!�\/ ��I�,�W��ƬƩMn���z�A?%�rKe���;AR�#'K5Ғ�=2&h	gX�5w>��h�LMaN�S���Cl\�z�Sݲ��<?��^ YũpNX���4�5��$��De���j�A�9Y�?���)Ȕ>6��KLFYJX���>(E�S�j8wE�k���$���4��FĴ����Wy")Ex�$ӴC���i���H+�OO:r�۷}YS	������m�$�ӳ�W��� R����?��Un��%�΀Bܺ�j��wHd3@����9�=�0FԐ�|�Y"�QD:-.A����}�;/KL�K���0@d9�R�?=hM9P�	b&A��ﳟ^�ϑKꌤ<������ ��ۗ}mmQ�M"��{�韗6�u�� �?zO:{�;�_�i$�b~�G7��Ԓ�����F��M�^��ᡯ������=�����i�p�G(a?�N����^���)!�f�;�N��a|��rKYN9k��y�*����l.��r�����c����S��c�}�m���֏�/C����8���}eׇ�)�k���(�%+�h�i���Q|ź�A��?��96����=�C����Y�t�|�yl��d`X^�yy�by2��,��v�
��D鑙J�@�Y�*�2>X�Fb��Q�;�v^K��/N�4ά�����ß�'����Q�ԩ��(}x��|m4�2j��W�O`�������rɅ������GP���W��sI�����W�Wftm�)�aw9܇�Q_��5
c�K�j˅�}}�Y����^��t����&6��J�~s& �+��G�~ُ�k��N`j��S1E���gr_h�T�v�-L���{��Θ;*��{|����5Ab���~�xp�����<ò��o��G;S��ac�5'J*��Jͤ��xrʓ^�a�	�Z_
9��5��c���� �Cb���p��k�e@�\<�2�Vj{Ehz=a���#!?�V� aV�݌��2��w��4{��/��D�c�_z���fa7嵽�vA�������?T2���7R��/Q������JL��	Przr��M�p�XSibg�p��}��=;R�����פl^�T��z��[�S]�d|mR�I���[T�燥V;�hCv�W �Ȥ���j�>�U�.+M9,��KS޾�;\���JM���hE��ta}8��e(}�j����xS铱B�:fՂM��́Y�E�u��'��dR�l>�x���{�f�j� )!@���@����~��F�^���4U��j����D�/�K��B3j)\+��l^ �⬩F=#2ܱX���p�8a�����_���G;����6��k;�+4��敒�N�s8X�G~*�evy�3�?� Xc�������Ƃ3h��sY�~�ʧ����o���ݫ�f���|w^�LUq?�X����О����)�̄��ԑ2D�gT��E�_��z#�h�
���"����ۉ5������Q�h�}��Ka2~{�`}��g�^�9�����}hiE~i%1�D��%�uSC�9����-�j��n�o�gd�a�lk�����+j��d�'�����S�ɰ��'򃨪7���>�ه�E�NO��75��I�!c.3f|}��X��>�d����-i�-��M�ox��(��T��0�}�(���&�/�
	�
��Eކ̧���	���w��l�αA����si���	Қ�a��K!�����bEp��Ty5�J�j�)�Ε7��g,�Z�r����v���� R�i�/ W{�|�wS���A��_lC��>����f��>�� ��7����1'�dD�>(���r(�
F�������c��~���A���	9惱B8��A��,�����0��s�M��P��q�L]�`�Y���׭1]!�x�2K�
���\�o�1�g[��$l[;O�b5�����d5�t�E��q��cj��D&(�Dٙ3S�U|Y���16_
�˗�[�ʐ~5��:w�x��l-kBG��������X��b�n��B�����X���a! ��B��׶��_��T��ά���5)���������dO���H|1c�ɶ�:�Ϛ&��ry�t��9�3�NR0����F~^_��h7:����Іx��������q�r
����ѪE*�0�0��g�1n�D��!/�vU�X�
H�'E���+����B@���n^���"&�'�u�c���������so�CTh��rZ�}nv$c E��(�(�?�V��_��G���x?<z��F�U;�>z٘�3=�.Ħ�Z�{�m�:�ގR)b�eJX�H`N�,��{��G�(ңk����@b|���&M�<�t��в�B�f��7e�D�2/̺]p֪ߴ�X��W����:�'�����v��V��MU�\Ԥj��}�y[5T��󨘻}]��㛅j��)�K����֤j�{��2���-h �ƴY+޶
�(�;����}�,��� 6��6N1���Fv_��6O]k���*�9Y��ܛ�l�=�%#I ���o���q9�fS��)�=���������w�0����dz=
�s>N�fB�n��ؕԾ�v��*��� ��,�M���!�;�_ݦ��ߚ_ fU�\�1��	��x͓a��Ж�͵!#П��1B�/�y�kqOb�ВL4o��3o
橥.~|�߾8��mVV�z�M?l�lh�1�֞�7�L�WY���13X�^G�x09U6r���ʦ8����	�����I�@�����	�H��	�,���@z�H��Y���/�75USu�T�>��=ב"���~KQ��B��\C�g~�޶���.��?� �"��7���{wif��7����0�g=qC1�g�Gޙ����۲e?�n�Ȩ�AX8 ���� �_u:���x��b5��������)�c���4jȓ?3A���`w��Y����!��Ӏ�L�n�q����\��EaY�ĸ�6�� �\�b>��(��c-�K�E�r�X>J}7�:>Q<m�_�"��z�����%���y��[����Ɏ���	S�K78B�x�A�+�8{�^ﳥ�&�(�������2�wF���j�LȺ��E�(˕��:��{D�3���C"	�:�d!zpto���D�_c�Ό�Q�BS����1e)G��`��L]��5B��e���؜Z��s�(�V��4�J��iڄ
Jd&��RRI��ĄZ)���2��wK�#w����$!�eI�ҏń��
n/���/��{�;�2i��\5ۜ(���W�7a+(�X\���#��do�2rb��^ra��Zq���p�nK�Tz�v}Zq]8jx5&rZ�8��B8��2�����Z��,��� �֗�i���0Z��aG�[��ǖN��S(.���_h:d��k�Q~lN}�./3O����7��/4�j�e�[9��Y[T���3�~]�s��9ڪ��_�>��CVR��c���/����h����P���.-D��pvASO�o�\!��S>�#3ۙT���S
33���5��?�~�X��T�zv����f�3�5�c[��Uxא48;%��rB�q�G�� !�m������u�/ ,E{C*)x�c�P0\>ߐ��UΣY��;�m<oؾY���Ek���#U:���7ybb'.��3���k�r�O�:~t�����kfdj��/�lg����������~!Z�{֍Tʷ`���3c�֧��D'�SO]��g����luP�Pt�����Ī%D���C�-�{Z&4��G�\6�������:������}oT������J�O�<E#�k�cږ�wTK�oP;>�hox1a2�<ե�_�$ �m���愦9H�m[��@$����� w�����1�:É3�>�8h~d_�b�hz��L�@�;u2�1α=�u�Agm\�z
b��"p�ƌ��p�� �����t��r�K��=҂�q��wA��p4(��F2�:�< �=!�	�Cꁇ5���3ef}�{��ġj4�8}q�_�P�IR����+$�$:-}���>t�C�
�ZT�:��Й��@�@����?�#|x�������,�Q�"��E��dG�
��vY
id4pd� kv��ʔ�����S�dV+�pp�-�MU�&�E[}�8�,k�`I�%h�O&#3�u�TKrC<��~<V�غB��Ja�������h5��T;��� ���L����tc7�Z����"ј�w�oV,�U�x5W��ћ-|$�Kx��?�}脁x#Ƒ\��E��-��I�*[xC*В>\���j	̖�<�> z\PΦ�y�?��4��?�a݅,���X��[�� ��3�:$��5�_ ��K����"ܬ����'�Ƙ}J��)r)��DL�/_PIb=mr囕�O�P�d�g�PF�Tk�	$��񲖡`�\�}����t�9�?�~*),=L�C��b�*[ʁ����w��A�;���	 �6W�*��N�V�M/+��c�䊟�҉C�zV���������s��2\�X���Ӿ���/�Jp��'��y�ofkn�K�^k�%}�@)K2�-��r4c���+  -�8繟�c_��kK�k�k�5� ��[]��e���%��	�3��D�'��|���|�,mKO�߬���AG�Ȓ�Iw�]S�U�d[����0^�\-�W��G��n�ٔ����MД����ϙ��z�Bu\�Ó�1Ǧҗ�bS�d[�2���%�=_��gaCs?�r�6Y;pSI3�,n%��1Մ�����"�g��X�w�/g6����{��������+�Rc��"U���F�<�a��{����OV� �1�$��Z�k�\�&�=(�BZ��+�_UPo��~������kf�O|L��L�9��������#�*���&�G�ޜl_�1�T,<�#6`����7>��`^I �i&ig�'�<o���m��?f3mz/���hNҤK�\�a��2y)�����B�ʈ��ٸ�y�1-�U���2X&t�B����*f��ק*J��%sy������8#�,_R	Gcv��\Td�C��r�U��MW4v �^-�4|hv��.��_'U(^�����s�D&���2�X�<s=�J�b�mEN'��ӡ���?�F+G�:��9"�tqI��?y������W��}c�)ʉT�)�~\���αK7:*�+��4	�R�x�	Lp�e�n>zLj�q��=ĲKy�K�3�H&D�G|�=���K��J����ُ���J�<ML,Nf%±�~拔]Cݞ��B4�O-=���J2?�@��\%1Q��PvrL�,.Q:��h���¿��_K�ѾĐ35�ba�v�X=��^zt����g?֛rw���?i��k�
sW	�6�h���՛��+��R�e���2�<)��(��]B�Zύ�O�3�ϗ+
Y�w��#�t���\�mp�s�qUoZKJ�.�L�������N��9�07#߄���[��)¿����@7X!�Y�%�|7�F��,�(2���`娔�~*��V��4
`◨C�C����:��kS���ROfr�A����MO��8�%��?��=;Ժ{�Pٴ�n���߃� �m;�tҿM���y�گ�X���W�(1���/���{�W����1�������
�8�+x�E�	�J&��-���� yw�x����B�5|���R�|�H-�@8_��k�|�2*Q�U���W��l>S��Y�K �EI
,���
����7��t& {�̽�#EKŘ�9|F�,�z��e�N2q�5w�P���E��Mcv�����{���-�혎��H��"�����{�
����ʄu3��@�u:����|�S�*씡4�
����o���)j,>�;���d�,�0�8´���5����G�9b�г�L�(=e�v'��M�w�A��Q���tS7�xId�C�5�Ԕ���R���9J�7�j�Q����hs�m��(��x����ݓw:},�Wh�p��^IYİƐ��MK��-���t�GΝ�m���P�%�c������s�Qذ\�B»vǅB�"FD 0��G"�͙kR�=�m��P����]���N
���:�5�J����Y�(���4@F��E-��ʽ0���G�K	�9a���C������MMW(�We�|�Yk��.�y��Aث���SG���>�-=g���-cf2���V������~�������y?	��g�3{uܖ�_ᰈ.��*>��~E��$�Th� ��\��k���fm���6{����ǧY�����dB�~0���dqx*�P�0�b�i��ʌ�X"d��Ӆ˅E\�Z�*��O4��4aA�;Ї�#�{7��҉m����-߃;�G�)#Ϗb ����U���\kߖ�i,�����*����NjWk�m�\:Tl屨��T��#q��-2Y����!�W%ʌ;$+p!as7�8$�Ֆ�YV[i���l��	� �+�a����^q2�D�O��О�Dۂ:`��/�R��8�Y��
LI�j|t��#����T��86w�9<�*B"L�I��4���Th�[��5�u&�߭M��at�ii�h�]?�l��t�R�#�7�+J4�ciC7���U�L�Z�����]��jO���iǱ4�)��0��j�}�-�KT�"�����}�?�W��^Pu/"��	..ic�s%�����@��+��dH�[�cѐL*J(�`e��p��R�S��';r@�!C�� <� m����^����dV�>�!�i�D�����£�*Ӈ�k]yh�8v\�\NIϺpz�'i�H�i(H{b���'!�p�;��@o��"/�sU6䫹#�~�+24���"h�����Us�a��J��&Y�H)V����6����eM���5R��RK��*�ˎ�˥�'�z������>q
/�!�,�u��\�C�4�":1���G�tѨT��<�f�_y�=�!���9�C��|����	�C����ǈxY
P�t����ɚ�K<|�8���6�����L�b��_!����@��0p�׸?��G!��D�B�F���uZ(���b'��1��� >h�u��.�Ej&���B?��_�~dԫ��O&\���q$"�6!�
�7~��;Y�N-�LL�1��l��?�:����p�R���Ty~<�W�dNţaVk�!ԅ�RAק��_�X�Ehj4dRD F���4}�3�bP�P[\F<RԄ����A{x��i��l���޲�D����?�q�J�"$������'*��.+�I���:O��ƻ�>
����-T^�_�-��x��?7\ w!�������yq��1{/�6��:��C�69�$Wf�ą�~vE��7���T+U��b�;P�V(���9�n$�� 	�U߻z1�6 9͖����R��d�wG-�ߢz�ֱ^W�C��*�R]�(���Y]說7׻�j��O�qL[Ȝ��!R6:P2��g��ш<�D�,�>T`�,��1kCx�0%T9���Y'����?�W��� 8b�u�R5gS|�u05暘ؓ�n��>/��Fn�Ys�Hx}E������y��qH�,$h��b<��ʒ�m����:�Y�po�twy��q��˜���կc�FZ}�B�����╬��%?��8S�p���[��rv�<-��D���Зa�L$� �?C�p���<Z˥(,D�C:s���g�b<t^lK�@�f-|6�8�Y��/��C�ؓv�맬�d*ђ^E�X"@c�D��|��i�t��}����ZpWMS����jWZ��������x��W���U1K�h��CB`b}o҃�׉�	FwD�EM�
��{V:�*��Y�mŤ`d(�}��+��tv�'�DnSk��� {�7�ؔ�4�a)�f�(6Wl��3�=Bb�nKj	R��%duzV!��K��/�Y�C'}:���$m8���64���R �PiLaD'f��j�A�J�]w̯|L�M�p�>�����������.Y��*�"OT`��a��+��"��c'�3�0�1�����ԜpN��8F=(����.����í,+ԕ�閂����P�
ކ�T�kOg�������PU~��= K�O۠ ��(��9(W
�ų�bW�����dׇ(���W�
ӥn�R���
��L%p`Q K��Gn���P��}ǩIG����Ht���$r�6*�Q��b�����VeTge���.�ni��;N�����r�����gP��<
� I߭�S��_ ��B6��6���Aq�����3Ɵ>�6G�/ w�ɲP�g����J[ZB�������O9E-$�}�@�BX��������u������9X���8A4' g��
�0��R{Kp"4c�wQ�J�\ݵ{ALM� �L����O��Ru�c������&��&4�řA���_��5��8��!��-�g��S��ҟ���t∝!���i�������*�7���q��(h�:\p@���bx�{hޕ�s���Z�
�W��3'�{K�� �~�)�dE*+���sQP{��8+�Q�
������� ��yB>��d���HS�r���KI��ܝ7��RA�|��$f���s��n�Tb~�0.��~$K��7}�c�6'��Q��Ww��B�'E�N�QUEYq�VŇ7:�x�h\Su�s3ȉ��֨b.0v�v�7wC[w�;}3!I��x�59RY�Y���9ػ�|��8;AA����J xZ7}��b�MG-|��.Ӭء�\V���t���鶺�z�@�<W��-J�0z��Lls�s5nJ_鴮܅�זW�~Ӌ��6nI�Y߇�ߘ��71v����n���y�-�`5�HKu	y���]e�H��]aK���Z����nݰ�!�`!��ՙ�p�D���n*��t��p�� ��j)����jUu���D'ߊ=� c��Y�T���}�?
��k}��|��!7(�i�y���)DO�f��Y�cx r�����J���N+��A���>��f��C�(������=B�@�B_�h�(�iT��D��`��db�a$>��ht栒&\�BI�ϪX���撎�� p){����#��$�0��'K�^c7<����p�8�y�5��0���*���Z�F�E��ߨ��А��2�'�>v}����w���w��1�F��*l�m��1���)d-ѩ*�<��ol[~�A���آ��G9Kΐ"A%�f��#��qq=��m��uumU�u&b��^�����g��]�p|��e��[r��q����;G��<v�39<�}|��1��q�MT����W�{���c�஺�cKw��G�Ķ� ����ef��Ж��u�=jm%}(\] ���h�mfN]�|�)E��N� ���NU'�5n����88��'�?�ru����'SZzD���8� �gU�@hT\SeE��q���C���T�r���9^=�~��,{�C��Ku:�<^+���_7^��	<>��y��	�xz0v[Uu૷A�_?%��l�2?-F;�]k�~�wY�Jq��S6G�iM���.S��_�R1�$�a
#��o�N$������g�7�W�ʧ���=)j�!Ă���O7o�+9܃?�HcK��f[^18�n&a��ot��_ʨ�hD)�q�d�U)S�)H���6�fL 	�"���u�����-Д	�l� ���������n�i��Ӏ��_��ϒ�d���Ǔ
�aLy�;�={򭢰l0,]�:��O��T�)@oa�t�9hf<��i�E[�s�n?q�8:�5;u<��"�	{�l��<D&1��i��	���
��+gA�� �)\_?�A��!�s���<����P/Yv��B���ɟ>��4��Q�l���s��ޗ�5��[# �\�%p���pй�*XH7� ���g��T��m#�1x���<���v$��rϽ���x0<���z�F'jkf�e^X��.*-�[��0����恸�J@���j8�c����r��֟��@��e.�4�\���S*EZK��ЇDV��K���fZ0����%�p�lr�޷�DW��S���ܰ�Ae�k�4�,������Xo��9~~��p�.H�=���xcA��D~�3AU4����!P� ��j�J��RH�Ԥ@�B�m�#q�4nϹ\�Qo�����{.@)��E��5�0���n-�����?�s�Kh�^��	�+|u*�*��5�*��s;���˕�
i������#@����re���Ѳ��z̃�c��
����ϵY�y�n�o��ɌRӘ�zz@����w�^w��-t�%�.P�ɑ0Q56]h00��P{�	��d*aF����ԝ_�����D�é?V�x��2sƊ�q�����n���v�%��Q�Z2|d� ���@�@�m�t*:���\���J�6+UUq�\�I8���>�G��J�#+?:j)B�X�^>��Q虲���K׀�ɗݢ� Tw��/�ջ|h�[��iWi�����Z�Ĕ��'߲�=��[���ϭ3��=�z<��8N��Y�+i'�n^!u�J��pa������F�C �6����(%���y[���`ν)M�hN���b,�T����[ScE�W��lPBO�F�7�9��zN���򃹬3���"�P����"z��x��)>i;Ԣ���,��1�����b�QRK�����Wy~�~X{�1v�g	�Ẁ���%�Ժ{��� Ȅ�3L�Z�<u@h#ϛ���~�`h��F[��ʞ4_9���I�M
���T�O����@1����¿�{��0�8
��h��f�5�
��kJz�F�@�����}��!�G�^��\���-|B��"������Jj"N�N29J������bP�O �;�~ ���T�!�Y�z�ʀ�ݠ�`�u���ޯw�C�:G��p��O�]��;Q�>um;D�睊onP>'4��RmU�Q��7��	��j��RIN����WX�E�!����'��}6w����� |_���e�w��"MJ����D!��c���e�;�^�elG���^�U�~D�(޼ L�\r�i���ܦ����t_	�H����ff�~9{F�6��4<r�ar�]C-��y�n˼5�z_�Kn����f�v�n��6�	% �v�����;�']����S�/z���~�Ũ�H�+�{cg�Y�g������T��<_"���:4��F3Dr��"=O����(Wԛ���R����c�.�A@?J�T~+`CL���XI�ݑ��} ��N�$l#�PqTaM,I͔�i���%t�q�0@�������3'�Dx ���#+(V��$��A�k�i(�3K��a�w��y�\84w3�q&�H�tܴ�e�"Psx���qz{Am�3ꬍ��ЩĬ�͋[��;3����U�v�ڢ	g��60�o?^ ����j]}|��T��]�ou2V���������\�ڋ_�j~@'oXG&*�n}xg�yӴ鄕��v^w��/ݞ��������kn*��$o�}�Ǖ������=��Wϋ���|A�����m�1���مϛ<;6'qB|X7���s�tٓ�K:�ǟT��,�(�#L�;�z���h�i�1�G���1Oܙ�4nu��o�J1��#��?�G����?����u��]|���:�&���O��x|��Y=�+*�s�HY�LyF!� ���SM���q
�uB���5��&?�����w�j��뻏��wΚ,=M-�];�#�Ga�2����(����6X�O��w7�m������COg$��OP��Z.)�{T<�s�]�O�}(1���!���5��P�R�qEV�B���]_������S�C"a�$G+���B1^�ڢ;��
?���
�?���>���������8bk����u�è�x�i2��n�_{�%�k�����R��#La�yFu��k�&�&5�����ʨ&t�~�G<�A1h*��'�-=�M��~���"�Ϻ��Ƭ�-�(�Ja6�����<�~��PV)� ܹ�Ŷaq�a�d��|��-�߀{3�����X��W��|�}1sK.�б-�g�SS�)��E��݊X�v�ڍ��@�֞��ԍ�/E3��}dq���[���|P�v�r�/������� ��ѭ�������`������Pݟ�x�q�2<\��IΛkӮYO���q��s
�N׮��\�i� ����)���,U���ws�S�R�l�祵�;��eu��M���5H��G�5�ZU҇m�ZIl�cըb(� 	rx�*��[��U��Q��8�	'z�Ѫ�?�8ĵ�2
����?���t
�,�.�3fJ�V~��G��?GVY!eױ���|2�C�.�l]A�TX��:3��ʶ��B�fv2�8�S(�(��8�b]Ӑ��)
 JH��Qb���K|�>){����l�$���(���bl^�����>�_��ș[�P򸲟d����+�<ia�\)��"�"4<����ܰ/Z��Ϯ�����z�����^ Sh{��^䙹��������Xcj���L�9)&cZ&{}�O����Y�d���MD���)�»���<���K�C�"�c_�d���m��e���O��4��v�e�RѠ�4�LW���JG��."���W������j� t�C(���2�Y�,ٓ~m�<-����)�ˁ�8 ��WӉeL��&�����q�߹�Y��d	����Ԗ�B�ȈV7>�Rҭ���q�ݼ�������݂��/ˉ����|���	�ˣ>�g<~y�&DQ��6O�bY��b%6�j�_���0�L�r�`^���g��e��b�La5B�ObX�wJ렮�������0kQ*Jt��f�8A-T���(�/�_=�D�����/^�R����k���4�3������^�s-U�8
�!��_�i��,5P�Lʕ�f�˒�T���B��{Vƴ���^�g�������6�����$ݎ�j�
��@р뚱p��u<�b���LQHMrZ6�#��qRuz�v7oK�! �"0P�� �&C!?����3�ܽ �ë�h����LRX��P�7��2_q±��bR-hIo���vw;�N���fȆ>z���!��'
�'���u/K��>� N{)y����	�='�Ҋ�C��Y� BFtש0��&����Y�R-B�2�GΧ�|��v$U�dT|��}�jl
^�ʯ��3�a(O�4�kzҫ�vi��-�N�ж�Tld�������/F9�++(��.h�X{����G�,d�ʮs��D>tX_}J�hnF�Y���C�tJ0�xdCT(%oi2�E��S�Ҥvɳ>UTT8�(T���,�IN
���Ƽ~��;�)\�&n�x��~U���.�N��n�_�=�s�Ԟ�%��3݋/҅×�dꨕ:^əhˊ�;$���͔Ь;��GLK���7_e���u֍��y^�1���Ѫ�n�g�O����{'��(�}b������3Q�W�P��]��z�hQ247B+�	Y�`���C�^|�ᡉ���/����%��($	�O�i�;pļ[u���d��e�Vr��oU[�s4z���T��� -�
U{ 2�X�^I%ۏv��I�3�u��@��2;���Ua�H�I�`-�b��_1�������Ssb��mv�	ķgN�SNY�#lpS� kA�a^vKk�MͿ&��?J�j���� ��Z�m(%�v!,�f;*�����y_A��_����Z�+x�����>}��j8Ϧለxxݱ��Ɯr+K�e�����T�Q쀂,��x�B۞�sY#]���e�Bv	>E�e~ef�I�X©f�Q��nlM���E��-�!3K5�����&��
���˘�G�d���x�FZM4ɿe�: ��B�'o��̊�xeRj���`4zq"6^j�� gm͒Y*$���)�hE��*���A�������xNU`5���N�"gX�Nr��N��0Q4��(�34oD�]���C8īd���MҠ���%���e
ka�,�O��fɕ���]xpJ�-�����pc%vR��u��"�+�r����]OҏmK�=Uf1E��u��Ol�����RKm��B��������s-�J�:!K��m����J�qy���"cF��G�(K���WЫGa����q��{��Ixa��U�ot"��0'g��;}��gbF��g�i3s�*90S^���=�_3[ה~��JŰ}�����~.t'<���'B�D��Q����B�k�_=��U�Эb8&�k��(���J�D$k���?@d`�S��1�M8a`Ef]�D��Eα�OI�;��
�%IW���ql3W�ݾ-��m̑��X����*���*�Tq;��|�f�n�_�
����2��˩����p��@����A�ѡ�#��n�p��1��G�U�X ��}ąl2�O�!z��fm��E��{%5�I�	��8��� uR)�z!)n�"���ҩ������u�^� 4��S���m~U	��H*=M��]u$�U{$m�<�4V��g�d�-R�|�@q�E�z���d>\;�2�%T�\��6Ү}��l�*\K�d��F%P(�Kp���\�p��i�BI �2��V�d��V9R"�Lz6P�
�Û������}が�bԟ��1����>��j�<�:�4ȑ��{Gs!�B�C��;c+ �ްIod������f������-����c%H��0�C�����v����z=t�M����F�RE�%;�����m�O��RÜ���K�����pCK�i�1�f�~ P�cM�Oz����x�$�q���%�b�0�; �����ѵ.u׿�m��O��.!�m|""��YN�r[�:VU0��UIh�׽�f����g�hL��G��|����2�]C�+ri
��*�o������㇥q�zv|ђ�O�n��r��]ݗ�>T��B$0�ny�V��\]�^�y�ڡ���x�<�k_��6�?�NL��45�.HM�
O�d�:�UNE�^c����H�3|�YN�L��b^����j��_�\V7�v����7��0Кj�_R��6�t��S�j����U���&Q<r.�Dg㈻E�,�o{ؘ��F� }���⃴�r���鏾߆�R�:�A��ݼτ�2Nhj�԰�pM��82/:h�U�����ab���T��[�$���$I9����iaA�AnmG7fmy�p5�l���(V�T���n�Ks�hlnߙ}�]?��l}m}:�z��M%<�e�ȫ�3�{<M�*fNf��8=ƼAa����%V�;���|O�dmز�@��ʦī8<N��	߉ p�I�pA��,9@����	��܆��h���]UK��C?��>9xr�q��MjL�\
�BJ�e;B*m�HI���/��w|�g&6{n��ݖbt��Y5��4�h>U9�$�n���l���uzv
h�G�oSp?�Ԧ�,�O,Lh8�̈�(�U�n����$��xx�-��b�y`�.?
�gNಾ��O�f"gx4��ګ3��T�����bo�xL�r��շ�llY#Z�)<9}�W���5�:��郞�k�ҕ�R
�B��xQ�y�Ǉ�Oe⁧/��M�O��ܩ��@��w�K��m,x-���#�ĝG��25���+,u|�Fo�H�%~�}Y~�,�]�EE�7��+�C��Q^Hy\=��E�aY��[&3 �:#B�S�2w0�b�S���OF�5=�8C&��Z�Ҝ���{�߾ѕ[�lWب#�J�)��(R��\2���W�/����-�|��K��3��YT	V@'*���6k�l=hK�w����¾wB��33�\�N���Z�@�X�g��&vI����mc=G��u�9,+p�$�V�wx��1K�+>�u#s��Tn|ӻ|CM4�����/�]�͈vL��VIT128�Q��|�R����*��;d�M�*n��TX�K@�'��8�Z�4sT��4�� d�x��b)E�I[�ݤQ�ѫk� ��JA=��\��������3+X�W�m���ٟLP;�e��]��)�c��J��]�(9��Uh�~�԰�$��'����8��8�H�v���X�!E�贽�ȁ�U	Kf׆f�����2_F��m�W���V��O0yT	�#r�7F��ծ>`ese
Qw�����CLt�,�T��L���Sg�]yw%������-t~3�k��%PLiGm��>�Ac��9��&��*]W����$;,Gݜ�+�u��2"�,J��&�/ ��o�]j=�Q�oX7�Mf�A
)PN����ě�v���ZS�
\�WX�Ʊ&^ՠ*tf��%��XW��󼁪��(*�P�VgpT"5�J$�ߓ��"텋�M�������.�6YQ8���?�k[�	O�r�#��TǱ���F��<ƭ%[����~��R51�ȦsG�MLG+���6Ȗ�К���{7�&2�UU}�,+)<�T�&�&
��'P��;�c�z	��Љ^�������?��Ct�Fk�i����7'iZ̧��n*�'������ڃ �!�5&��v]�)����gH �,�"7h!/?���"�/�G�c���T�~�!ұ]>���5n��g��FQ	�Dc�=kɗ��ވ"������0��L���Rq�95q��su�ӆ�	�HƁnI��-*�$�N�\�%Rn���--Y��i�}=*�b\U�����\+�oa]�C��ܥ9j�Ɉ�j���?��B. �'��ӝי&�,MڳrUZ��`�����usa�u����i�Y��:tJ��˓�U�H���}:�O�6�}m��.酻��,����B��CV2�4ߘz���T��j��RU���ڐꎬ�-a��uv��[;s�[�ɡQ�e����+*̹�Gc�e��Dg�Q���GJy��9�[ SYu*>#��˹U��Xx�A�ֆGc\%\�'8��K��X1|�����*�`rYS��� ��]�D��'�����@�i����D*������Ӳ<',�Iָ�}�d�p-��}�%߮+�>�R�M\�Y��ua�k���%�G_��r|���_�d�T���}Fc���c/i4%��w�p�78X��A�J���d�7��ܻ�ٸ�be�9Fia���-�a#*'7b��l`7|�t%�j-5?(�i�m�C��1,.�N׵�y�����"� ��~����M�k��׀��?J���,��a��%��+q�8'�Z�l�^�_�i���A�P9������g.��c���v��/��)������y��rr%�l��M�Ι�B�zz��}9�95��N��s{p�i�\-�qi(�H�}���������K4t�(<���N>į�,l�y襎�9rɗll���Py�%�!:�U�ꭝ>��nE�+3�-�ӓ����1TǬ�@���],S��&�Vت[����,j]ȶ5��|�b;�y�LF{��&��_e�u���
�k;���������h�#�HQ�$�)��T?�p1��ʙ���k�r��&�xE�-�N���&.]������n�>��n��gc1�Qe�?�$��qr&S��MÖ`���ESq>b�� لݦk�y� ��΀>���)�	w#��ĻbT�53��7笃���m�9�3�7>P�F8�zz�H/$Hl(�A�b�`Ib�T��~�t����
A�4vu�n����Q}��\�paUv�ob�2v�(Ud�Bq;:��`A�[lA�����
�������@3o�u�}�j�;�4z׶J�֦�,�wO�g��0��r�| ֹ��Ɨe	T���\:X�o�ME�%Y���ؤXa�`��eS�Üi�����t���S/�@��@�����6���.���U�n���!�Ds&��i����f�d��S��[y�j*f9J���\�TKBޓ'���:77Y�>�s$(�TL!x�]|�y�䭨E�N�dE�^�9��=@ݜ_���z|�gÕ�φ{��镁�Y&��Fǒ �t��(�x�)�۬ Պ���&���x��Ow�GS4��ٽ;��#�%LL��,E�f�d���P�W�o>�(r�!fB�$><?������5�u�F��pgs}��.��]C��j�5��Z��V�e[���6YF#.q#��c���kK:py����b��d�����tK��uO��pM6+��s�LM�`���5&=�\>�[4@|��̗p�n���Ý���JB��ơK�?F�'��n�����8�2sK[���T�̋���.�tO��.^i�@� L:��k2�j��oC�yG~���7w�ݱ��H����]���X=�-��F����q%I��Yk-�����3KC>1C<��\ޮ?�u;PfR�IV�G�*�?>��}��R�>��������w�2��N ו��S/�I����
n��LO�� ���L����mo\Yg�ܴ�rٖ}T�����|W�庅��c*�ւ�\�r65��5Q�_g�DaY ����5Z�B�r�ɒH�쳮��P��חG	,���J�t�i�i�f^�x��M{��R�����W���/ �G�k��<G9`�c9�Ɂ����Y��Ĝ,^2_�
X��fܹ�%��l�Y���1�xͅ�!/��3��IF�}���l�L���W r�F%.��J�5;����5�А��l�>d��KrK��n)��y �CSy˚` ��  ���WjAL���ť�BcY��Zt[��=���a֔-ւm8�*�ZwW#�g����<ge<�� �':���C~h�C�A͟$�$8�{s�?� ��?�g;C��f�-Ӣ�(�*�ը�Aj�n�1�r'qk� 	�ED�{�g�yP.Q�{���[Т��s��g��_�\5��| g&Ç��3�z�/��T��ʬ���S�5��|z��Ӫ
 q+���Vx��8���+׬�����&��.�+�A�J���b��}������T�����ԃ�3������s�#fƼy���j��AmU(�k�����[aoC{��qp���˗�r	5��c?��7��yC�F�%��G\�_q�"�RI�*����%�-5��� ���˳�?澪-���v$��@p�%�@pw��\������%�tГ�\���ۺ��<�U������5$�wWWͦ�*�v��a��F�����p�1/4�W����'�3�l��� n�/��
U,�}0�6�Rc���T�
-��X�2,��'g�(	�y~��P�*�#p�9J�N1�;>_��ȣ�4�`����4���ni�6��e`~u��l5rI�g�8��$��(�F�r��2����`�Hn-�d��#�d��2�T����'��B�GO�E�j;�}��+��ӍZ6�+��͂�L�	B�p'l�q!���H�:�d���z����[NC��:5U�����y���o8A��F(�x\��pO3a49�Bp����q�#��L<��C��v��@{���99w�C��Ֆ[z�l�>b
i �{��=G�aF��u+C��1���(^����ď�6��p%E�R��\G�?��楀鶇�9��vc����/������Υ~��&�Q�ʽ�A�oך��ݟ9-����Q�P��R������F�N�U�d���	��X���J���5��k�ދPf@�T~��ԧ��y����*ƴX�+�y\� ���^@}���*A���*����f	c�>X���L��d�+g��)*EmJ��z��������"��$�����h՚�H��L��T�D����aȂ�SlD.�׳@{Gs�+������3|Q���Cziz�0h�K] ����3p/��G�Ky�qv}K�n�-\����
���Z�
����>Oc���[����mx��rU��R�o��]�()+T��������	0Cx`�=�����va*�>C�נ;׿ޘ��6o%�U�����4w9|�gV��
���|�KY��C��/NvL�
 ��ʨ�"��4�����k��O5�R����|�\'5|�lR��U�Zf�k��z�aĠ�}� �X)=��tT��7bv�JI�c���t��*>��m��8��3�q��+����!�Ah����SrEO��$�![6�˜JQ'3�Svܸ�
@�?׊���2+1<�z}l6B(�
�f+�)�Kl詆��%����nj��st�T}A5r��e��A��z��~<wlJ>q���iX�B	��pGW;��I8-�ǌM��h>�u�A��s������Rm�c<Z�`��q�ڜ|U�	a?w�)Z�L�Ԯ��j�Q��� 䤱Lz��@y�R�m?}p�.���h�����(JSҊ]�K��TF�f��`ϒ��n[�Hx,��������S����+ж�s����n�SO��y(�p��+����8�&WV���de��HXL�Fp�H47��t�p@�N����1�t,(4n.���m��	�nߐ9���]|�]�q����b��Y�lM�r�2]R��k��9�|V�*_�8t�+�K���8���|#��{|�v�쵹$��e����o�����$P��!�魖KO�H�	�-M�_!@�\��:��^�7/�ĻpG��v��B�V�(�vum�Bqw�����Ψq�l�U\���m��8��>��T3�K���p��l��C�4�2��;����P���0T2�U`�vG՟��	Mgi�r�l<��@� ӌG�@��aue��U(uTU(c����'ӏ�z1c�z�ZJL_h�iYFGw�k�Bi198����Dwи�Or��.iJ�ф�?���*�ے��R�>�OS��H]��R�Γ"������^�T��ʐ4���*�Bd,fuJm��w�}3�������f�fC���w��~p��/������]�֫�sk�?�YI
w(K���]>�j=�'�aS:���$�#�V�~�.u��W;�}�pݹ��gW�Ë�ߎ.�%�Fpn��)��*y}m6'����� ���T����0dw�0) +���'@=\W�z`n�`'nI16z�����c@.r,\@��N��k�����}��f��U����8@�UJ��v� �O�8�8�G|8h�r/�X�\���Ϸ4��[�O/b�}:��:�>�v��4�v	 �k��I����}K�&UR�Ƈ+T���4�G���#�EP��34��++Ri�=��q9
�I�C���g���{�/zaE�i����\9��Jzh>�G1p�ٍ�i��𢱛�6v�Y��E��ɥ�Nk�ɸ3�vQ�Cz�r���K5�C��<���tU�[R��"!��ऎ��0��x��}L;Y֖R�nW:�b;"/�ۿp�Y���(V9�#�0��s�KМ���=�0�1^���r]b���yO(����,:�2e���C�q}E�|z�N����;�V��aXpU(�C[�G����T7z;_9�ʷ@�,\'��,Jyy�R��v0֊O|�$�H�%���+uJ��������w�Gp+���{�����M;}����
P~���Ƽ6�_���d{��N�̩�4�l �E'ߒ	�7�/^~-N�3jV�7��՝��c��v���"S��1�tY��D{��l=�a��䵎�-���Tk�/KH�|D�N�f?�OYkkB��sT�W(n��"�h�\�БH�3+��R�e��H�Z�]���S��&?#G��T"�Gy��3����K 	�
M�~�>�T�W�f��a�.��l�v���؇D�~21�S�T���<$�@�a~ܽ_'�� v,�9�ڏ�R�zn�`�d�tL�T)3�f(�?�v�G&�r�,��d_�s�"��L�)O�-O�Y��:Q _�3�U����=�n�y x��^�~�/����/�����6�tV3ޢ��\��4^�G�H� C7]o=z1��[?���8�D�����NX�NW��o8�`�03�:� %�4S̲ıg�-hr���)2E��7)�ҙ~�*�h�@O2/)��Hp�-���:E~|T?" �������j��p���x�]������Qx2Y�X�t�����\<4��4�"o�{98��6t�#6+�y�2�Uś�p{1>���K�(I}M=B�Jn���hs�㳀Ԡ��K�lѻ(>�����S���"�)<���utC���뱾ƕ����8쉚
X�^��R�rW"�x�G��S+Ey��Q�>^#��x��dI�Ӟ���0�닉1���n�^�	�nؗ�OBU�VeR��-�59B��I�PD�dX�x�yi��.@Cٮa���F`��$��,�qtpy�A�	EIC^e�M-H�|�9��_��O����2����Щ�C*�D۵p�t	��߫��(1�����&lF�<?�4��A�(W���[�U��B��z��?U؃)�X���-(\����P����(I��\���:[ !Z�x���.���$��&Q���ņ?�Z���e�Z:R��߲�p�vͭD�|Vz"�f@������5��l�/� H�h86�F�P+����.������x RA�8D��E��xf	���n�	��/�~(�	�3�Fns֞���g���Ŏ @  )���L�m���/��S�
Xӊ25��a?Ἦ�D�,���z��[)A?��5뇰�Cj'swH�\|��mp�'ӓ���/���M�W�c��yS��+�}��ʡ���v�Mi�%j���xd��:)�4��������Χ�Z+#��dv�rb�
�o p7o�ی!N����2��>{��;Gmʨtuj>�������<icMOy����@���p����9V���]�_���YldF����m��$�a e�-�j��4ѐ勠�1���Ñ��BfO����}���Y3�]��r�����@�+����|du��wJx���#�����T%X�^W���_זɮ6���#W˯�*��a%�5t6��=-'ò5?�"(&�cr=�^٬�=,{��b"$�$"���lr��2i�M�ٟ�~~ֈ
�'�K0mQV��z��o�נ[���c��{h{C=�`��Ֆq��>��H�3�vM�=x�`Z�Y��Kw�^y�yn>���W����I$��G��"�ĕ��S����A�	���̹��ݥ�x#۱�\�AL=7b�G9�8e��cB�q��Y#�3�]�8� <^���Cn^\�+�b�
[ {Ȋ���k�xx�R��Z)Q�~q'4:�,\֛kh#�H%X\�`����K��~�X5<�Y���E�ٺß�{��u�_�:܍0?�|�aý?H%�b����[��g�E�'|#��O��hǙ(
��i����얝}Ś�o`�m���N�Z�ӲuII��ؤĲ����\/�#�9���@��{��	����3L�!�FϹ?��r�v"�^�-Rk�C7D�-r8���X"-���)F*h�\\V��R���w��k��,���mEic,hܟ;�HT���,�R���̼�
�(�D�8��
(˶����N�yea�X_�U�zY�m�sS9*�$��%o��΢����Ρ�<?צ���`�ã��
�ow��.�Df��OY�溔o荞���(����L~���m*?�2d�4�o�s�2y2�صz�=��B)���t՟6��)�ΰ+�q83X� �'	pw�R����`��c�$k/���:�bC�����Y!��L�������5T��&��D�hG�rS$��
��l�yS�"v;sg�o����Y���� �t��h�9� ��Q��Ca;�X8��D����a�Rl*��AA'w�l��\�������G��ރm��ㇴ%�x� w&�8}�&o��Ȏ�s�
YG�=���Wi��f���k'�ĔQ<C�,�dC&LM�C�C��V^�˸'��Y�ɟQ��6&�3���Ps�8>�]t�P�m�:��8G<L��ԚA6�tdDD�`̧��R��y�K�|R&��l�. ?}�?��ͫ�k��L*P�!����QUU#/����-�4uѷ N0!>H�n2_�K���4�yZMHR�p1_�#NԵ��t�H.k��R�̇e	�7o���F?J���S`�Ri�;k��M�L���z����:�����^���9	;H�"�137}�uR�Yʗ7X�ԅj�ZUܰ�{X��96B���N��a�ݞ��5.4c07�pm2^]�^��hQgBc!DԻ�F�+_@c���7�Mv$}4r�
K��Ϙ�nZ�
�xKO�"J�8j�T�.;�"ޒ/�?ᲠR��Ezv��T�>z��L��Akn���]ts5�ī��H�FP*0�eM����\ {�%�F2�r�`���g;��?	�M�uɲ�1qJ��L��aK �R����H��X���u4��ݬd(85�X⋊}u=��������2�1�ܐ1*�n����R�~��:�!3AR��7�\�")���T�{a��U�M��P�MMA�W�	��	P��o!�Vp��_�,���]():��]>D%�)��X�c̄�zU���"a4�������;�qH����+ �̳L�&Z7�}U���y߿��#,_�G��v�R�ۜ�Yq��Z�������v�qe�1�P�lQcn��ho�o����u��
��m��T��`�7Z��l}#㯟�̰�hT�ցћ�%��D�]��VQ:]t���E�w�D��6I"_h#�?��p~�s-�mٰ��r��+H|->�kv�-43��8�E��E��9E���6S�κ�y��]��] �5f�0W�������*�vѧ���#�cTz���YM��)�1�%���i��4�L����$©W���4+�9��CO�㗏�WG���0�c��%�����X5��k]*�|��!��t2~���"r��	��|#��*ԗ��}�2bQE��}J�~�ʣ˫�T��bF̶3��z�|��?���8�1��&�v[)�]P�R��Y:c8[�-�{����CM�r�8�\�� ��c�u���-ǭ���,؉c)�3�k�8�KL[�+��~]�~�pč֧Qe U_�|��ոpNTv#Q�'����P<��T��d��P/�;����%�H���L�$�W�w�@�c�N��?��龤@�<�� �s�Pmݒ�Þ�RE(b�5�_����P��|�$��H���}S��c��8�O�)�Q�2������{�������Uq�x=�=VU
�f�%�|������fc0,@������ ~]��Wb�����Sğ�<�R,ЀO��҂^S���������Ĥ2�6N����'��N���v�6"�Q����k�eJ����Qދ: UR���K"{|[ż �A�nн��NQ�[��J�@]b%�> �*aT<����.=3t>K���`�S/�Z��%���#��P�-�C�̹�#n7�R�F�p�pM�pF�����xj���3�	Tɂ�D�V�q�$TK�V�^x��᳉Gu�$�=X�@�~�>- �K��:��������+����Mz����j	6����m�.2Dz��B��	n/D���NƘ�.���2�G9�3�@<1�zI��.���%�y׳���P{��$�_R��3�d���r ���m��ݏ�uod1�}_�jh_�eO��K��s�P�E_������,*��7᠖�Rh�6�`hg���1�ԝ��`��O��Fkg|��.���R+�ڒ!u��B�=�X��>�!6��R\���?�$d��v�d;���
����`"u:���N1��3���~dk93�Gh�[ ��|�Z��22�W�<J�H�o�5�8'C�N�M$���@0�܃����U6�~����:�)���IUؓ����ߋ��S$nfy�1h�|M������/��J2ؤ��E�)p9�`���S�� �
f9�@�W�{�ո}җ7�d1�����g;� �4�V�6W����[7���OZ��d�:+ݾu�Ш���~��b�>�[�]i��u�3*���	G�2^�ʂ� �ۜod�%Ա�N�C��XM�0q��#x��A�D�)'�^sU��ڏ���I�r)l����GR��]�ӊ=V4�{�'!���,h<=�����.�ԯ`G��$u�.�Q^����tE�e�%Lx����"��y�H����F����E��d0�ߕU�I`y��}V _�b�frQ���½���	�~�}�W��w(��>��M�����R��0���,�+��J�rxk�%νQL�õ{�Mf؜	��"J~���6ε�nXӊ}�y�Q͢3�������J��Kj|8�eΖzL�+@�+l6�u�R6�Q�k�cS<�}"[�pP���tXk�=�2@#"|�vB˛Z{�t:�۸���|�I&&�˺�x��8�>T��������i7��%�ۯ'�ID$$�����ij�����i�̻(�n\n�H z�ן����g��� ^I����?z8~�q�0���ɧ��C�*�0�P�����p�+�<n�m����̖A��.���)@�ʼ�j-�
��+I|L���R������+@U!vw���̉�EJ��B�o/Sl0O�ɲt�V�c(�������|e��5�|R�5@á�Uv������ޕ"��M��4R�`]�J�f�z�{�tj�h�R�p��·?�S����ױFs���gwV����D��{��x�58<��LƔM<�}�X�[�q2�]{ϸo
�O�s����Dz�i-U?g(Y�P���)DU���^�/k��
@k��`,�
�:�U�l[t�皙R_{�f�vюR�DъuLw�K�;б������[��`	A1H�;�F�E2�Ix�9�q;�iz�h��ļ�Z2_!!�' �=[]}(�������K��a��)>p��>�,�oU�H�H�i�B�)�����ѭɑm��췱�K�-���Uwv�ߓ��	t�*��|S��eelhb�5�X��Y�ͷ���3]��+��ҁ�l�(����y듺A�و/�W`Ćv���`Q^^i�9jh1E�\�� �D�Aw�� ��d��;�Y��}6�X�Y��T	?=�(����pJ�^({M����f3q)�mɋ/S����+�|����� bo���9�!�J����V��Z�VA���b��ƒ�}�L]�h3;��8ei�r��2}��_�֦i�#��G�0fÎ�͑�ȷ66���:ٜ��ј�̤ͪ�X���O�c�2�j�����b5ͭ8}}WI�S\�Z���}��<Z"��*�5��$-�}%:�'6*��&*{Uչ`SS�j/kչ,���_&��ӳ?�Z�Q#Q4����|'���?mB�ղ��רV�~`Iڸe�ɨ�讶��J���W�31��S䕽5`��,�X��I��W���ɾ��x8�U�$�:��L���N�}S�@+�U$�Y([K����Vt�frG���М F--b�B�':6��
���Q�jn�Ue�7�kc������  �^n(jʤ��]C�~0��J�G3�c!{ܑ���T��+��H���ِ0ؙ�3b+C!)oJd(��񅘡2#���/�<�i�ޣ\��7���2�
�Hy�b�&Ȝ���M����+G�0�*�R� Sa'&�{)O+,~J;Zc�w2�;A=Rj)G�S�N�<�*g5��_ۄ�,�\�;ٲB��)~]/�d\b����s�C闢����[hۢ�T���xW(-�g�-ɗ�.jj�z�n u� �JWCz�Gx�+�K)���'���3�6�ƶ���Ѡ�u���x�&��ý�xy���B�w���x�����R��+���z?��e�~']���#F������R��ߒBij>upS�Uh��b�W������J,ֶ,�b�F���hi������+�tus�J����i�#:A���d�i}f/���A�z��#F7j� �.N2/Y�4͸B�2U;�K��Ո/CWPn7��8��"(nJ�^�48Tx���>�.�xn���)�S�bQ��7�?Y�h�)�5L�6�򟣟;�U*
�55h^���4	r�|�!�%���Ś���cD]���n)�:�b4Z�3>6E<B��К��l=���;z�.F�s��
��L�HJE�A_|�}+R����^�<�^@����R�̀	ؖ�C�u�n�R��Xq�`Nw���6���3�k-��N���Q�lj�{N\��N(Т
5{��eUS�Ԕ��f��\c 2��m���Z��jن?��x�-��؋!]j::JE;����ru�w�G!���υ���n�C���	2�||-f7��F� Xa1�<�"�/����f���0U���o>�ٚ�[�hxuz��'Xر\? 8Mi��R
�2����m��Y�T��R:�6_�DOn(���~
*$���|����UF�=��R�^t����|~ �?ZKB�,���]�	�x͕��W��UQ�����+J��12�m��r2ԍR{����dv�4����s�8p�ėkv�kj��_�N��n� yy=�ϖ�X��8�n�Q/���}*��$�x)	�������]��oBC��^?p�e4M�~�w3����kru�4;�+f�"�I��X�6��+CR���Q�L���y����"���|���/P}��:j��]�x�h����򥟽oQT��n��\�j����O�8���VXµQ������'���m�k��mc�[��X0�W:�MEB�@8�2��)8�[(sUE	��Қq�'׎�/z}�_~CW�G�4#EnU�Ҳ�7â��;?�U��C�m1C��������오�>�f�)[�N����p�˃w|q	���Į�����k����>���Z�UޡYdf�H������B��)g3��:��Ө���,J����(� gr*U&�nԱ)Q	&�	����Q�)�闛`N3�*�+-M>R0��f��g��ц�N�ߺ����,���M��J�?�WW�1��=˭�Z�T��tk(��)3��*��c�t�)���@O�[�.�])@���6�}����]��]3�SW�۟�O{��hM@̈́5�_�a:TB� q65/V�n��%�j���Ij�P�E�fj�5_���|C�����tj���������''������n�'j�<�W]\ckdW[����2� ଳ%s7�ç�l[�O�i-�oi��YЌQ(�ҡ�R��f�4ߥN���n��������5x_*����ݷsy�6F$2����d]���F!ŲW�����5�vG�-�bG�����Ÿ�&�I�(�����4��b#�^MzV�ӿd�����z�����Rt��T3�s�h�mg�v��M�
7�'�j���l.I����.���S������lR��;��nMyŻ3��r9���% 4k(E�.�~�x��K�	$�-U����ip:V��.�Э�v�X�����)jOV�ꩵ�bP��}�0�h�Ms��^9>j}�"��� ��PZ��o)&��r80�S �յ6~yy4�K���	�N��'4�@�s��6L���g�Yq���������W}����G.4���YZ�c��y�d:Q0pm�:<`�՟/��C�k�����y��C�����r�'��)V�	,C�+��l����I�M�eq���@���T�1�&�c�x��~�BHHi�/ RP��8��1���sG���w36�M�˽Y5�:GH�f�TV�d�5C������/�^�:�-�y�\��7�k�\<zc��I1ƕ@N!CJ2��Y诀����i��w$X�?#�	
c��5�X����2��(Aن�S%'��O�njT�:A����H�BA!����~��C��i ��̙��7f�H��R{��E��
kF_�d��񬯂��s�6�y����Ǹ�[Rե�tY�!�\��\� ��k<�|�1~� v&rQ�E�7q�l2T��)��[IF�;_Ԉ�Ϯᮻ��F����H�ht��T�����VV��Y&������1�� ��o�j)��!�a�9��-7)��s�:I�c�J�p�ة� ��0���W@z��X�}{���A�ɠT����67S�EO�����/	��c�����h�������6����ZU�����u��wQ��cH\�ݸ��ǰڮ\�h����&�.�(����g;�l��o��eԘǹ9pY��{f����#�E7?㫿�w��M�v<Ty���[� >øT�������{��V����w��-k������ު]2LC[���!�"��?k�G��<?V7����Ȃh4Pn����E"�qe{���(S�tILv�aD��뭙 ��I��oi���}m��>�!��ð[��Yw8��k�+A� K1�H�&�H���F9qG���z�mg�f��y|qDᮽ�\&?�yv�T��yF�dE/��i����h.{��z��we��D��,�9M��_�2��|���çƨĿ���ˑ�r��Tjk�|� �#�:��Y���s �/ɹ�J ��Z�m�n��{x�bM�733_`y�I�[5��� �;xp����*g���R����Jߤ�z��Y(q�et���_��
x��.�]9��x+��9��Z�)�����L1s�X[�Y��η��\-�I�=6��-���'��g��l��4J�TI���o��DO|���P�cb�D���v3;�yƻN�h��Jz�q�el�5<µ8�����L&mh��V�Ϣ������9h�l+�Ԅ�H0�.�*�����Ap���F���KL�+���3�������Q_�E��Q�#f���������3,�W��+:�j�֢rbH�r�X����o���g�ِ���1�����>����G��z6�෋�����+����Wz(5^E��F/�(җ5��u�E,Uu� ���5�Hؑ܏(
��{��J��k��ڳ��3��<��˷eo�����ꓬ���P��~O�P s���У�\�U�K��:�ޭ���2gxqC�X�r`�Gk��_ʇ,od��nP��f��N�q�e�R6Ӂ��d��5%�V~���x��4;��f�x�a�Kc5�)��y§�ce=����%�ޘ7ъ_���ZL�	b�\�̢Xh>����U����V�Bۜo:z�Ϣ��1|��b���N�=viur��5�W���+��W��e�`*�Ԯ�k��B�x��?VD�0Tgۑ�QZF���J��R�-�='��:M]���i�n.	x�,�N�
&d���+l_c�#$���u�^��ϐ��!��v�뽣-Mk������w
V�%��FN���J�HG����ؿ�qw[_ݩ�Y�ůV�/+�hݗ��������iH��?�$�Tw��m��w���N�!��EyR;���a0�q���exc��h�T�z��6��/��q[3Y��"Iu�«:����P�,(Y+�k+�5����� 56�&�-�6�˨�fdN�J�
�v�M����Br�.��d.����;q��K��������.�ˣ3��&�V�1r��(��O��lI�.'`��ЊQ����.:��=�&�2��
��'� u˯��]��V� O��h�z���NCG� �b�w��2�ʰ�K_d�·���
�<ӽY_�)C(�yD�K�eAx�NQ��ʻ9�p�(��e�u�I;+ȅ!V&Y��"�f��C�Q��,d"�	G�X�1�Y���Ί���imA��H���Ţ�8���&O|�3�n���>-�C�Y>��[�~^~}+�����G5��6W۵��7��e,�K�ŧ�Ǣ�J&1�r�����,�äa*g���"��x\K�C3��E}2)-�((|\��<�ZI�s��L�B�֎/�xO�Y�oS�w\�t��xL��.jb�F�Ǎ"GP�.?� ō�i�J�aP�u����ڹd��L6/�ך�����l�c�:�[�i��A�/M�?�*ǐu5%�|^S�'�$�Lg����加O��?в �H�:ѯ���a�sz�%~���;h*�|��e!�o&�XR�Qb�[�P��-PԈ���m�bT�8uV=���~}��3�׃��a����`�xA4�lT�*��c��;�r����17�q���U�PE�ph4������t��ص��W���K�1��%{T"�wJޅ?=8�L�2��n5O��{����ۡ!։Ē�������P����/6+�FT��3X[�i��sPdq~n�m
{O��lR�@+��$h� �i�j[b�0�%�0RQ*��fG����ȴ7�8���hy`�避����&r��]���i��aIg��c�ttt�H_�DXc�AA�tT>V@ZG[��c�����]��CO)�_���K�
9'1�7���%P�C-�f��"+�x��ޅ3�HD�lϴQ���/�?[er�U恲�)��*���R�VZҭVqk���<��^V9I��9}Pu_�1���CK\�1����$55l��G�
�U����^�����
�����W�B�3b���d�	��yA���_s�C o<y�����x��g�Eo(��ß;xr��DA��޻^�g��ԯ����Ԩ�
���\[�/[O+k�/a_����3m}t�l�^U�O�㺌-j��`Mjb��͠IT"\�N�3�2s�(��<ٰ�{��q�9�(L�2��UD��%��̗nI��/��eBA9=��!Fݥ'��P�,��z�o��A�XŀZ���=��a��N'���+�0���0���4��o����I4��}��M-���V�Lzb�VY�uS�Ѱ�|Ɍ������������lm���L�;���]d@HQV᷺,<MEa���������G(���[`=��2{"�o��� e<K�4,��ۛ�+����"�$V��iJ��j�Tx��ߕ�j�M[��W|a�����Z�r����H�OhFT�C�Y�*�g��ZO�W�\G�@2H�E����	�����p�
�*����l��F!�����p����^��$�oZk'��++��o��R�hѼ��{说͢�6��\/G��o�d��������mc Ƕ�vnU�~#�,��-�/���a�����_6l��2�x8,2���N"G�4�y�Ye��6�+rˋ�͜�N����2��[�i�&+��FH�/@JDK����K�}Mu�!:��=���@���!�i�ͬ+ej�}q�_E�k�ecx��k���%�X����o�L�����V5����=li��Ƭ��}��I��\m��0�"՚ ���@_��'���A��Q��Ƹ��J�B�dz�X'�\TX�t�������� t=����:>��};dmrZ$�/ȫ�$��9�;N���T��'���p����y���rW���%E\@�$Hh��ȿJWVZ(�D�0Y�C�(��*���u�E���
���* �*@��v/���K����H��fzL*��=����i�pŭ#:�"x7���0:8�0#d��=��-Y�$����-��˲a�%��()d�B��N���K��9�s�J�E9���r.�${�R����Z�,���Y�Sʞ\������t=�0��޸ўګ���7�HI\�<�p�P�
D�Sޤ�3�$�-��!��􄪫~�,��N���ؔ˥�ɷBR]D�$,��xd�S��ĤQ�fN?Y|��.�{;�q�nO80�g��r�M9�g�#������g��v�@.��B!�^�{m%B�9�����q�
m(��s3#�O|�tU�g;x��u鬇�_�ik)Rz���Ʊ�'�<��
(�o(���9�T�1��5A��=j_�Msm��oziM�"���q'qdL�VN�d�ɒ/M��{��FՔ>1 ޞ��h�T1�G�K���[��sv�z��݆�U�mLC��"@���c�}�^���X�̄7b^s_\^08?23�hVǉ�py| ��P�-��ں�g�����jt�v��M"z�l�����T�'�Y�=I�$�v$�+9�}&Zh�U�ӭTV��E�H���;�ט���"��ۅ�p}VPS�ͦ~�V����6��ˬ���v�c���P�['Q��M�ì&*�֛@�W�t�;^{Cۥ Gcx�rM����YX����_�����lB�	�W��8��Tr-j��' xͻ�F_P���uO^:�A�\V�}��>�V��zQw�����k������9d���w��l��n�0�M���i�`/CxC@���u�xy&�^�o3����v|(\<耣�G�������q�Qh�O�_������%��Yb���_$'�
���rl>�����_�m,nk|���T���:[(���)���:�����ٍp6B�`�'�4�pL���yQ����!֕2oAY��A���iڍ�������b��t-QCB /<
��q%�"�P�KA���w�JM�j_Mis��D���B����{Լ!������h<;�wҔ���B ��72d)��
7^�gAm��z�����l�,Ab��q��4�?$�J1�ɨA������<�o+�O�E�:t|��"�~���}�W�s�S���C$�FRR��&'}֤9L��`u-5¢j�\a,�,���v�"�ˈa�)�:�K�QO�D��a�|vvѦ��}��V��=�f�ա������%��AȑR|�Ф���Y4ޏ�'G�Oy�0[vt���q\aӂ�����qos:[����K_�����r��NkRZ�)3Z���5�4��0Be�G/2�aJ d�.���5e �Oj���[��k���+3���<B�O�9S�)����y��;�SD(_K���y��^:���s�B̪7�͌�lt�(��<+�4���P�]ʗ�u����X\�`��T�h�Y���)ե�_������$�=ʱ�0<��`�����ݧ�S{������¹�.��Î�yX�`5��V��~}P�@��|W��!���ڧ;ӈ�ި����>�Jc��H.�c�OK�zE�_=��[�/���E�?�\��Ǐ���}R�B9��߉j�l�y�����]��Zh��>����riM�,J��V$�����9:�A�s&�l|;��0�A�J�Oc?Sa	��[�Ԑ#)�k���b���P{`��n?�64)�O$-��dYoܬ<�ٻ-N�Ȧ�����j��3Mp��7a`~���p��ʋv��	����= 8���I\=G����E��q��M9bӘ�%�w�-�,���'\��.��X������69{y�$��7�>F�i��%�Za���,v7V�ix�
-���w6weF�����_��&a7�U�v>z?I}��I�x���� ٖW~Wj���hw?&w�k��\m�ԓS��V��a��;�@y�߃�����~G���q��n�@{�؟�;�b������z���:V�O��
E_�)��ټ薳�$��A�g��@,l]�Q%9%9�R
����l���K#���J7KH��]ҩ �%�� ���!!-݈t,����>���>_f��;��9sD"�4y��#���[����ؼX�t�����`�R繞j�9�;I�{�(O��Z�h�,z���.�D+6���h�z�+g���	��e�	����� �3��G��w�w����GI2h���KW3& �Z�@�+�7�m'��b	o]c�+��B
�� Ӱx���jѾS���q]PPJ��� ^�>���{8��3}yxd�X�����f=���d�[�ư[����=fuS��CW�IQ�	���x�W���{G�K<����q�)�'�n�������Ҽ`WOV+�	�C��&Utq�K�:�=���#o�Pޗ3�ў7��˸�l��ME��&ȜYS�7T2��/| �a"���-^7�@�Q�1�s���}�
���岬�
�A��#�b�lG�gqܙNjޞ�$�������_-!LA1���n�aq{Rzz��fJ`<B�������{�M�fS���῀x�*!^��{�}q[��}�}�5�!�U�8���3I1�к��y���R��E0���)I9��-CB�	ǡ�\;��П��T����V��n<�2��2g��7(���?˃�B����9���]p�o�x���F�(�u�H��A7��Q覺��V-}�=J͓v����"��`�f�7Ct��b�:���w������)#@{��ݹ�-6�gz�8nITV�/*R`,���6><���0a�D�/Z�4����^�x��0�r�1�w�(Lr{�M��jR攆��v�G���rDT��cW���"87�oaK�Zl��c`�΄UUNpn/�v�H
���������"�#�?�J�[�ʉ]����0�9s-��%04�Զy�Y�c�����p~j$�o�����D���+U#h��Ezsj��z�4�%�� ���+�J���kІ�1�C���q�z<���ݷ1�zE���WM]�"��X����(ŉ��������?�p]�o�"��O:�[�t�iޖ"������l�V
������\��D��^t&$���2�h�Fu��rY�j�۰�HI$O���;�V&���10	p�jr��Q�[w2t�����zBxҙ+e��z��+C��Sr����%���_�z �7wǢ�������?Zm��T��4������@�Ø*���l)e��}��H4YK����_(�"`�����@s�JA��qR�7������1V+x�l��K��]��ʶ����2`ט���]�����:�a'�#�-K�ii�8�镚ݧ���Ҽ�!ip�=��aV����O:�KN����+�++������T���)�3?�!��A�d֪D�1�8�Ǥ�����	�W��&���k�@Tw�Pw�q	J��U�?��FK��c�[������#�^�#�o��<{%��v�!��2��%�L�ρP�
���پ�$��z/��#0������xlu�>[��4ɞ��ڲ��sN�F��@�k��-ݧ)�q]s�̨���.��s��V��j�70,*�Bd�tmd���K�u���w�8Q�	���+I=���ߛ��#��+9N�/Y�z���$_u����鎪��#]���J��8=�>h~���܍������ t��a	�H$�L#0����8�7��D������^��{eg�N�;c��}=�~=�s ��	�ԩ 5NA=;��O{�P1K&��#��q�.^4��b>�|h4�h�U�#��� om5.SDKy�<�_�aO�$Հ����l�޼j�[m���#~v�O��k�����_r˓�QB����m�\�_�:-� �+RU�	�'�Cq[I�V�vc����)i��ǃ�#�g2}+Ttv)F���P�rw�,s�`���A�/u*�U&��&$���f���֞�{�����',0Bo�n�1��&K�'�@R<N �]B�6B��gysbÄ�d��r��K�W�6_�K�L���K�$x؎#G\�p�^���I�j|�v ��Eb��j��<����c�U��,��Q��r�`CS{�GH�0��.��p����g�Z��ZHd/*�n�o�ا��U�Yr[�TJ��<���c}�Gq�������Yŭ�@0;�!�*-Q�Y�jx��ک�RjX���rN��Ou;P[���Q�����)�sXW(�[�H/��jj���Oy%9�\<���}�U�h���V2��3j���,8���~��^-^{TsOt��_�b��h��$�p�RI���	��}�L��՝�  �*���&<���-忧�F6���O��Z���%%�%������o����؎����B�.�)@��Nlq�.aA������5�����;�<�]���Ԯ����sh��ѯ��?�&�ܴ�{FE �H��
�\!Cv7F�}nΒ'7��Wh}�$��k���-z��ۗJU�2�.*�a%j� �J�3݀:9Ոc��Q���֯9�ּ�$�\��eŵR�"\�^���@Gۛ����"|qq�H.�����$j�v	�y���o�2uxS�\�*s�؃+��T9�
 �f���D����ɲ���6
��"NfEjp����"����&,��yG5����n�U�GG�z3bL^zC�Gg��,,�嘍��3��<��D-��W�̢�ձT�/��4��$��o~�ݳ��dd��2��pup���}�h�oߤ��ɰ���~w�J���R�Z�R��������� �s��-5��"��ck#��˝xJZ��U��?kG��vK>��E�+�ʩ3|8�<е�n����^vhZ3�(����X���X��,��k"?-?P�mhp�I+Ć����i>�R��_���=�0����^�!�w�Ed�do9�6%�s�27�xUΟ9�f�i���C�H}��Ws��e��h/���C�ŗ�oz�1�~-�Zi���_�E��wj ��o�Je�Ѭۙع>>Iн˶�]�i�m�Z�و�~8B>�x?��N�~�'���+$k2�_B�:�8��9J�A2��ΡSs>�qn#}�N������b�,Z1�!-�f�Ƶ��Qix���\�>v*���F���"q��|E/u�l�[S�!aW/��S��E�����d��B�:m:42�Y6��NV9���W��`�=�?��d�®���4s ��o�9|�/��,D�X�1��C��a�n.y�p���e��귊N���S��7���2Ѿ�ٞ��L7?�qAW��9������ i��ѿ�%6�C�17���^������u6�m�,�^�:Y��\G��ו���w5��U���H�`��Q�=�[���Y��%�v���*Nz��X+�߇��#U9�c������=Ri�����S�U��C�}�Lٴ�W�A�~n�5�� �U��B��{%��w��\$�Q��DZ�ęT�,������ z��ƕ�䚄W��	�S�e����fA��F7�����I�^7�6�?2ݿ�ʣ?�[x$u7��7����I���'s�Y˓Ud��y"��o>5�1���o(�tVTT�̽��Ǔ��}h�7�{+��=�%�����j�U\%\L/�U�`e8�
�=xf�SSge{��ݵ�d����AT�r�f��t�n��+{E�zV*Ul�2̋��6���-/���&���_1��OW��<.��NQI��Q�W	�O���`�>�l�4���5���rea�
��Z��Z38� [[M�s2�[��;k�H(=Sp���b��aDEW�}!ۥ����Y|i~s� ������`4� �\ᆂ������X�y���s3��[ZY�V�Ƚ�ۼ� �cA�;��nV�*������ڵ�}p4)v��l��#���l��d�*��>4��ȧ�7��R�(.!�#J��\cƍ���f�ƍ�/Y��	���~��`��_@Ac�f��G�
V�b1:^�!�T�]�V������B��#��J�3=�Fl�3E�ӿ��<[��]�q���&��C�8�L�
�?���v�͖���|�OgK�hQ*�ú��jHމ~X'�B�.�Z$I�B�h�"��J��}��S�ʟ{�U��)'Ä�` ��f�.8\��̋e�U
2!� ���"4{V��I�\W7_��PHV�H3�HD_���C��x�-ט���Z��+!�����ͷ^Ph#~�Dj[����P<��|�s?L��X�K&����&�uł$Ă�����#�P��*=3�e�	��E�??ޫ�6Jȍ���|Aj||k�,*����<9˽�6���r��Rp��Z�
����Kē66K�������W��,W�#�.�P��
���;j�3!H%�Bn΄e�����jL��E`y���Bj�q��v?7���J���7��Յ�1>@N��.q��F$���*����>U�RO��6����Y������H�/�뮮�~�o7��`m�����|�⚟���[I���(�B0������V ��7���|e�{X�i�q��hU& d�����"�*R �)"X��EA��5�Q�;�s�N��*q����ʴ���\���J��+�h�� q�2y��]
U�p'�6玞��g��{c$�B�2P��_ kO�{�ØN꽾QYJY�n�ϡ)4����,��G�����w`���Y�������Y�A�}��ݯi�i�+���a�����1؀�IU]�qQ�,�f&����zj��÷���)���%�Bĕ���@�x��)�U�O�{�A�-�J�!�P��~�e����L֨�Mb�.��f���r8����ċ��C~}���{f�����?㖎8C���M`nǬ�Yb�'�a���CP��������k�k�����i���{�t^ u��t=�A��=���)���&� ���3�/�$UY��%�#4͈x�=m�'#I��x)M���w`������Q���Ɨ��~�[%��g��ttI�#N� _�ߠD$���m�+�y(U���P�Ɠ�dďi�O��8=a�����ǎ�3���ǟ_7�nԩ�bM�	�Pa�e���h��r*!@26�V��k��B��5R�[j��?H����m�����t�R�(�y��1�Z��az�b�{�UD;w%�f���"+�1��5te B�ɬ���@³���H*ǅq|,����*���I�R=~�En�	*��Y�B�����!n�L��S���,�_�z�J�ð�_5�6�za����˖�O�O���"��,�j�}@?PLS5-/j+�J.��#r�/��:�om��,�I�UvP�΋��BmףM��!`]��o��k^��j�l�o�?��IO��Lk����'q����1�r���|�n�]��BΧ�����o�hNu���U�x��iJ��W*0J
�J�距ϲ߁��h
�� B\]q �.(������uZ~$�$��]�����<�|n<�J����$ʎx�I�x���94o�C��#S�;$2�׋0��
D�6���B�n�i��_!��y=+3�C��_ �_�eཱི�C�a~���3�8�r����8L���H�3s����Y3O�<O?��V��߸#Fa�����Wش�/ ̛��-slp�H>P��Xo��D%KGY����<o�CAX�+�7��61v����ǟ��_c2#c��w����N���~/�9�)��w�N�Q�=�����0��"%��)��zn�\
�7�!;��uC
wҼ�m��J��~���ho|��2v8���-�4S�&ct��D"ܙ���N�8�8΀����KL��{��nBd㴿g��#�CZM�F���x���G�M������6�e���߆5�2����r������M���r�D����	�#�P	h���3��G�|���@j	m�	b�٦;��e1�$�O����g~K���F�p��ɨD�)޸�s/�cg�D�K�	1���Ի�÷>�,П�_^(�̈́9e<��eI7J)`y2 ������qv�<�� ������4K���fa~�䃺�mP�1��b�.���MF��-ޑjϑ�`Ah�4���F��װ]G�J�%*��c��G��o�"W�n�����ٔZi�ЊKVƪi�����H{�����y���g�)w��=-cj���C��1���J5v�ٲ'����$�P���� ��m��� dVP�p��y�z�-�����IrU�֕��8�����Bx˪���@+�El�pwMb�~h���T��n�UV�SW�q�le��ʦ�˦6�����Ħ����
��d!dIB���>4��L����q�|�j�4��/p�����aRLdC7k�F�m�ކ�:�Ն���⩑kMʬ6��QA�(?�R���j�x�D*()�;|ٞ������O-���7>����2ID��ʐ�������-&�����@7��BA��fO�J\f#J��UUe!���,�l�?YV<-��__�4L�
��ϸ��������_�k��W'/�� 	a�����\ͱ:���㥍�E�s�7 �o���W�6���4�a5t�������(ȫa���߀~i�;J� ��W�bBN���
�
�\Y-���s��+�m�42�Y�,���X��&P�C�r8B�6aO�jHJ�Li�[?C�
*�3X5��&.׃ճSE�e44���GK]A:n*q���P��L3@�7��V ���~�w�3�l���4�X��Q��\��a.��ӡ)�5�'~�>�L��m��d'S&�G����}r�H� ϰF���9��wwܩ��S@�'�����h`���i#�,��<W�q�U^w0!XYi/�G��<YT$�bsV��D �7=߯Юz˲��ȗx��p�~�Z��䇷�&�~�jG�Ji��[@'�$�	R���#Vi�|c�+IG2f��κ��a5�E��[݂h_ �6���[���1��s���l-�8���v~���w��1�vB��>�4_ �D�>�?��׉�q*�|��#\�|b���h{/,,���N�*�c��SA_De�ĳl �
��i�~�����0C�Uh���-�[L�W�l�F��!-�����лY](W^~R*:iEt���&���>��A��_)�K��G��ws?դU�_7T4 ���n�{O7�������yĲɍ��O���h���\`�v����^ ��@���.�R߅�H5C&t�@Z,��ш5�/n��|�v�����<��U���~��e0�t���繾fܬ_�示|�#���=���ǩ�DlG%��J�&Ӣ�����wd�����O���½#k|�srD����ƞt��V�S�b�r&��!G�̶wHj��̱�'��RH)K����#C�+'5�Q޷�<��5��r|}���*wz�z����$��&���X
�^��zz[�.�$\�y��jK�yq�vudT]]<O1;:p���1����ڠ'm؇suu�C��|��lQ��I��h~Qߪ�aX�5XN���f��c!'�M���#���T�G����쿸ʩ�Ri�N�����~M
��	�6�W��2ʴx���F��\��"�\Y網�By��އ[N��)+�37�4��F��z�ij�;�h_2+�6��s��3����S`"<<���7��Vd����K�gr�kt"����� ��C������-�2�1�q��Tm�?��c'� m�1D̀~I��Z��L����y�c�#��>�5�����4�Ԓ�P*�ô�0q�QCdJ��(�xC���y7[���A���>J��&� �@�����F�wTU��g�*�����g� 	�MmFӃ����z����ˡ���t�x^�?g�`.ӑ-�j�χ��;%��o���O~�h;#33�)b�ZVf�e�y��.߁~�L=4�upL�M4�ɪ����S�?�à%ɥ���V�r���z��\�4�衚��?��"�����eQ��"n�v/+�ʺ��O�F�khe|�j�1��,����w���h�)�M/ A��O����9ݻ����"�w�?Nd��LT� $I�^{���\(�Ο���QB� Q�)_*�A|ep��}�o�"g�0��wK�ZA�#��������O���}	�U������TEy����Qߚ�P>�?�R�X�7o)�j�ᯈo��1��~\�+�h��P�Ӫ�x��fz�ַ�	f/E�@��+t��e�Ms�|�(�t��I$�Ҿ�P�0�zk��Bg=��$��Ƈ��)�69s��4}��'s�J�%��?���	's�m����ؿ�{�/�����������`�-�"�L_�r\�`geMK'�/hT�t��k�o��)Β��op�x� ����g˷�Q9˖
��f��A�{�wg3�^�� 8*~�I�|�J��|�o����5�}#��eD�� z=��C�)
�q���a�s�ȝybAꁾCa{�ts�"�ܶ�0�i})L,_�ֆ���͸B��A�7��tk4c�ք���(Sd�mY�sܼm!N����3~(�8||�/T
	�'�7����������Z�MO6�NC�Ҧ�~v���P(>����,��c�L3��6a��!��Av`#ۣ/O�9��N\H��M//u���<�o�=�g<�J�TN��پ��V⋋�ڈ5+�� k��I�;�3*���?~���U�>ж9'�R�]�Q���d}/[�{��Y~k�t�Ɓ�ɜ������l[\VEsE�)[1w��6�C�����qC	����'����x2NC� :\�~�j��,��	�#Z៉#��+>���޻�U�5Y�c��X���@����>g iQ��޼ D�jw��BF8����L�[g��7��Z/
���z���w�T9M���煰����`�M2̋s�Y�|r�^ ��Z�fh�c
��+����Y�����e_}
�p�\~�2	^�+�Ԙy�Q��_@�s�^��S���%�p������y���FR
͙nop]r)R��x��:	���k�S�*[�@{��E��Є�?����B�~Ħ�s�+j���Z�^�Q��'�DSe��
��b��	-M�K;3j����v�,w~`���W�e@jr���}P#h�-ȕ�I̜Ӑ����
8�V3��_��َ�F����0z<{P��g�(!�}6�sJR���@ۼ�=^�f���"��!�؄��^��Ҩ�88�O�*��龨WF�\9�2N#Q̒��|nИc����=�C嬈�V�zVUW߂�b'$�- Z�����(Ȯj-�q���|"���OQ]	����	�� ���Z��3��R����!�<na�Q89d��5ߪ8~�<\C�م[P2a�wd]2Z<n��j9УDo9֩УOL�h��d0�����h�R�۠̉�gP�O�'��v���4Z<� $����{t
*�, �}O4I���A��bP���Qtж�f�2&���#	�K5:��>KCt�8Q�/oOu�l$�q�C��JK�-�`�ȟi~�װqķ����%A�ּ���K�_���"e���=T�7���R��z��!��dL�D�8z}z�]A�@
� ���&��̴u%��2��J���&b�wi늂sL�=��#�X�\"C��}��в����Y�_ �u�XgY��^��y!���qv>U�����Eϖ\q�k۪ۀ����~�T�^�
��x��o�H����Г$��kic�󭄱Z�=aw&�𭉭�1�:��������A�����l��u}G��GG��H퐠�Q�W{�j����DE�n��;�{�T���U�G��1��m+�A�����S
��+��.������V��s:ہ�CũN�0��i+R�����w��cc�5]�����By8��V7P,����u�ر��,���vMH�ߠ�Nė���p&+b.� !�@�
L�VU�?$��H�̷��PB�h�����=\����do���H�}��(Jx0v�;غB��Րd%GU�^��GK����"�n ����e��F�Uΰ�߫g��B�F�@H�JfXzG[���b?OY���/VD���b���Z�E�\Cd���>��op+�CU���wm>�X������} �����B�Eߓ�i�p�
1H�j,��Ҽ-�wY���� ���?�#���㗋�|8�<IL�ڣR� ��<lT�CJ�^ Mw������kH*�������C�-l6�yC_:gx��m�C��w�Z�U����#���p���E~c�50eY��-ƶ��'��'A2z��Y�׌r̶������ݴ5�;yZ����gg�OI#W� �a�}o��S�d���EL%�%9�*U��ōz��d�茚ݺ����e���(��߬�s�r��
1� nH���7�5�2�����ɿ�{v����m].����Z�B�%�|�L�$�i�cִ�z�M�g:�w�Z�I�R���ԩ� �-].9�]3(����I03���V�P�^�w�7�7�lBW(��H��H��PVO��44�$��y�L��@�tz5��|�{�j �j\R��	�F�(е��Y~�RV��}��:���HK�����⭼���L+ƅ������[���Bwiѻ�y�$�Ԏ=���o���Dld� �%���t���l�U,[����өFy�sI��T�x$)���KX=����v��:�L�P�t��H�@������D�$��� �Ya�{+�NU�=�¯識��S����<�<<��l�$�-��42x[�$���ud�&b6�^�&@�~;��&yӘ���ͼPT��W��9&I*��	ٝ,m�d<�����S����>��M�rX����{�nc�5M��4�:�����B?�3=WP�@��@~ڇ�/����(w^�f����H��%���eܧ�.�ۊH���r�6R0�V��B�Z��̑r�������zr��o�m� L�e/������P]��V��{���|�x���}��$����-�ާo��[�HΕh�HߓdB1�T�!��f�Lk��Lp9�0lի����)d��5�m��@�2BV)L�d��x1[��u�p�Z���2���ުѸn�A$� �����$�4g�4��	�~���l�`֌�D�(~�P��Z��V�>��N�U0�w{1IUr��^�`>��g�}?I�Z�nt��s�!`Cgy��aq�\6�s7�A&�6lc=C������� �8��\��K���\n��b���\[_ ��>U:�Z���=�T�O~�{;�I��|���h�Xלs����Bc�S#k��nc��y����v��"8��%�`C���K1�<�`����.h��W��-�Z��b(b�^��^�FKw�����서���k&EҖ�Ŗ嚥�PSQ�AQ\��%	����fJ��
�"�\Z�����܄�`tI+q��z#��umZy�8�����TӼ�5��)欎LރU��Z������mtf6���7#N;�M���C$��/z���r����J%�4"�솦��Ü��U8�d�n�>?���e���� ���� 1@�Z}�s`��e&~\�?��PeԆEz�3���C�_>�R�糓��qPV��BJ�/e�E�Y*�aihmJ}@�cS��!�)j�%�W�㯑[���^���s$ s�.���He��u�����~������_�-5 �������컱U�YpTI�����w�E��#�Rf��2�������f/��x5��82�ڦ��������{�8�!Itfʴ���e'�tI���oe�� ��'+c�ش�@�2W��o�������G�V���̈́��1�0	�*�a�����|Ŕ���l�V��ϋ��m�����B̳��':�33_��mB\v;C�<�^��u�6n�`CaJ~f2��jm�?�%���;aO�*x������|PgS��9��EX����:Q���,��
��\����#a�Ĩb;�!�âe�E�����>Z޸�v��4������.�3�����&�˾��-��"fۥ0T~��;�?mB�p��� U�������S��&7�
/��w_�g6��sI��M)��ǹ5$4th
��2�^��_*0G��{=\$�RO�_7��B���DE�.��,v���1���ʎ)���~��4,LI�Xb���+��~F. � �"��8�l��m_dE{A��	���n����,�˃�l7T�����)ӿ>!\ՙ��c�c�x����G`�y����6��-jp�N��M:�2�N�ep �����>w�)Uh�}��!<��ե׶ ���8��瓭�X�(����������7�*��V;�ɤ^����4�2���|d�����#	_W�� ��CTr6T�T�b 
"EL�]��a[�t�n���q��
�W���{�v�{��pȺt,���뜾��Q��#Tf)��r�&MR�NҬ���?N�4!_�kD�(k
]�A_����oZ���(L�x�lv?��A�P��Og��0[ C ��h�9�#�
yV:+o��6Vۚ���a�Hz
���?��F���g�`�UDR��4������NhR;m�r�a)�y-eV��]B$�!ߓ��6$tU9TK���1�D��+�&��+RG�>{��R�?3�`���)���b_��	|��"-�U� f��]6�*s܍�D��SH)�(�*�����H�ί�4��5��#�B�ǈ�U��2�b�������wo�}��e��V�E�l���ɪ��T��a���'R�s���1�ټQ�6lA��RCe���Jm`�ǣŵ��]���g�`*o9ۙ��MS�%Lc$+��|��X��5>o!�r��_?�d{H�Nà��,Uh�1�.��_s��+P�˜��y��?�OU�i�|��/p���2=[5/�_I?��)�:�����e.g����)P_=�1n�pچV�(D;SH7�&<��Z��}>;-�}t�U�˺[fO|���Ag��U٢':��T1����zM4MM�M\^��xVL�pnv�D��p��a�w����폕X�+��@J��NUhm{�"�di�D�5���
z�F��K9>\r	�̊�¡N=ӒNq��j�p�`�NtN�Ӌd���)K���0V�S�/TR�8�@>�2N-��g��-+�?_h?1�7 �d�g� ��Exg+��U^�W?��R����9����|$腐'��Se%��"�s>}��LƐzOj�L�]�P���p�K��+.���@v�CT���0@���Y!��6<���Q��p�p ��!�É�+�MNu��
	�=�P�Ae�IwKm�#�ɀ��gZaIgV}������?EQqo��+VaUh���b�8% ��L%�I̧�پ�\o�\Z��%cL5 �m5���u�`<��P���ǚ��%����8�Dyz��nocy{Tn�a�S�v%��K�R�8x���7��P�W;lh9jYI���O�!���/v�����,�bUz^�R�7���'��j���q�3P�u��(���i�d�~�X�f�1��Q��=B�ǯ���x��+�����g�=2���߹��I�g`Ͻo�v�<v;��7$u��7-eL�0?��Rm�,��=R^���4}�ʟ
��V["�/%*�~-m�.^���Q徙��O[���D�Uˑ�Ԓ�o�s:�!�+�E�&*�ķ�b���XJ�6���àɂ��xnV*����$h�	��G�Ky�:	��H=�O��� P8���%V�7�Y���V�*g��m)�z
�̍dLjs�nEڎ���6`|#Kb��0 �l�fȓ�/�_YxM��L�M)��`��~�0�x��tf(�_���b ��ҫ�ߒ!�*l�+$�S��w��G˝�߶��J�\�;c55f�g��$����>v|��v���^]��ѵ]�J�|H�c���}�ƸUA�v4([ow�� K�z�{���]yK��-�3,$�1~�m@:�	�9�Ѳ_w�w�_�*e�W�I&g��sDo�~��������#�������PX�L��.}��А������e�O뢩2o}�*e��5���؀<��w�JH� �zE?�d�G¹���Ѿ~ꜥZ����%f����4|+Q��j�M�s��_�}�7��,?}p�P˩9-�i,�~�����Z2pK�L�_�ַ�Ry�yw����퀘|yl.�h<�Kq��Y���Ԃ����y��?��A p�B��WB��}�e��|��6#$�(p$юf�nB%���dz�F9�o����C��/j`�ryX���RY�`J#��[C�j��*�u�Dؘ!��\��uK��ӪM���A_��I��9]�A�xa�[���z!_��,�gD�&����,�$
]�ـ9�y�e��(���^� �O�\�e(�g=d j*D>�(E��;������yjO��|]	p��(�����I�����wܾ �6�ޚ�z�Efl(R�8D4f��pu�d�@�$�!qDj���� 5��v�+iIN����`j	Vn���&��rs���ʚ�Փ�;����T���X���n��s+�Q�X��D�v-˸4�e���eo��^TQ��s�
��1YLKCōo�!c�X��Մ�P�Sdd����Q�R�A~��Ҭ-b 2{�x)��R����
�Oe�]T��&ʇY�P����1z�9�@R��>�5_]Ʀ�o�M�v�q&8e��u�6�c��#��5qR:j��i'*�r"�|�X�V��;q��ǀVŰ��,��:z��&֟`Cx���D�l��*��:�<���O�?
��>��2��(EU����+���v�z*^^:,����z�k+��b�Qq���so�Ǖ|��?�Z��̣oKB{z��-��c���p���� s��p��k��Y-b�f{ӽ�U  ����q���4VVD�k�V����E.0Q= ۓ�Hs�&�o���܍�g-"�^��?�8#�R�+�j�t�Yx��2�
7eq���}M�l+r�/�ת;��b�;R��҅&]>��=�V��g���q��M[�8@��O\bu��<�@cA�0czs��~/Y��%I��i���3�Ր�6�n�`����I��w��b��3�#)[�0�b@��	d���7�j�p�����Gu�
i�>Pk]��ly*;�Y�������R��Z�&�Mm97��Ո��]3��.�h)
@�6f$�l�1��[���o�B��s�ƪ�L)U�,cgg���,2ؿ�p����H��}�prBb�s����-�F�d'�Ԃj�4�7PĖs��C���Rk�Z�Bf_�eyT'�&T�C[���/ ���#qèS�>5R�%��]�֥�\r��*u���2�Bcٶ��2��pC=f+v�턋B�Fps� ������t�r�xx�E��}|~RF�k�|lq�霐[��G��U&]W�I� �4��w��V�<ST�9����B�y�U������c�?�Zi�V�/ ]\Ew���g�B�����th�T�9�����
ULG���k�/Uv�vW���v���X���ɷ$�U����=�������r�b��R��:��8NW�_Pm���U��놢�X#u������_4_����[�sfq�
B�ʿS���u��/� M�b|!:N����2��J~����)CA?��M���c�,�T7/�:�t��|bw�+d��T�2�Ѳ�Tz��+(]!��|-}z�P��<.kEO=�:U�N�~R�͞����b[� (��^ 桊�FiQ�A��/ �G�_��I��XF�)'��]���j\F����L�css�Yy�&&FB�
$��L,t�e}���Neh��8�C����s@��f��=�:6ڲT�i>�yV-�r�XQd��
:��L(����G�Ux�8n"(�srp�Z��vZ�t�j�Uq<�uU��Ȅ5�� ����g���荴�~V����a˓��t���uԆh�3(F%��g����}X=Q��ULT�l�y�q�a$yb9�II@۸�crv���ˠ������������W݃G�K>[*�G�O%�9��^�_J�)���xDX����Է�[3d�E`��u.8"�YL�G������@��O���)!w�G�m��~v��?،��v�Z��mi�'����ۖT(���ߡ>M[j�%/w��Ma꒪���EW�;���a�ۆ��:�4yV���L�2I�Z�����G��3W��`n⢤�jb��tU=:��CH'�}ؘW}�@���rEX�}��������Tl�Ҽ����uX"T�m��s*������#�<��z���z'j�U�K!��;��%�wї �kH�eW'z�V����W�.���y�����9׹��>��|�̙A:�������U�&i�S$���ޱ�y_6�m`�dt'��I{����^o�Zv���m5!�b�O�y��anTd��e��~�>����d���3Mx�iJ��Њ�`F��ym9�n��9~��y�K_�4���|%aF�%���3�)p�Q&L�x�v���K�/k�([�=��E�t{=bĤ�]c���{�����,ᇑ�� �X9����O˚����vb���L��-؊}�����1�f#�~�*<,;�"� �U �P�sګ�3�~�Р�9=�,���N^\~Lͫ��pQ2��`(%�*�C�L"�#��Ō�tx����Y�"v-MĀ?���+o��=9C��X�B% d���>��D,�&	E������T9�q�o�^�zӊK*Ò���$�͗י�v"=)�ʺ f^I���&͢`�k*� ��=ꇕJ�WN�ߵ`��=���(�V4+H��`W�b�w5q!�?3F�g�y6�S��������#��Й�
`�7�2yt��`Y˳ߣ����+c�m/3����C�`5�샌I=1ҾGZ���=qa �y3�T��9�&XIC٪�1�n�r/F$��ui}a�@ �A'�����d�G�>[ ��曣��pP�"!��(`՞Ĺ7�\Ҽ�����N]�'i��˿��j`��O�b�)}��?�ϴ�'��5�~�߈N��^����q�>%�� �} �����s1�	�EW.���N�kR^J��)^�R\�k㜯�*-��I�bxR'e��[��rr9�<'�^*? ��YH��a�^�$,a�5�zp.L���p�x{Z;:��v]�+�@���,W��
9��YN�<V�����P�qv��;��OX6������yt{�,�}�l6�,�/H1V�s�#�6s.�Q�]�a$�?+| �ȇ�= �1q�I~�@HZ��=�}� �<�m	�P���t7/�	V11��1f��JuD�l�9H[1��RP,O!Vz8w�V�6Ū��W�)�g�����Ň>j1ڧʨ��`�Ml>�T�}#B�����c�-�>%�b8u�od�O^��֣�X��
𷜐1JWe8��k�=��~W��x�}�|�$$TN��U:|�� �g�w>Pp��P�U��M����I�u�oM���<k~�n���ͷZ�P���I&rdpy����Ԝ��ڀ3��8��~q�z�[��5� ���u\�A�{R���H��V���kW{����;P4m��3�P��U^��t����o��`��y�ɛ��-�7�%��?�d��V-h�}21���=>�"� h3�1~<�mK����iSXY�"3��3<�2��=�i/�@�)�q�aT!�ZF<�?O��m�R��`ԙ)�x�	�Y }y|;�i�Qd
[��I�bD	���j��M@�򠰼�aܓ$�����?AD��C�z|ۖ��@j�]�z��{��C|����pƸ`����<���N�SȦ�)	�3ݒb�D_�kJ���I�������o�L�f�"íagxf��V��»�F�� BzVŢ�5�{E���xkN6�4	T�c�WtE��i���lA�<�;%q�7,��Ѱ�/{uy�x1�,0��Y�'�ԋ��Ӟ��]�^�N�o��ʷ�� Tl�o��HZW*��
�R�<:t!�s,�� 
�L���}�H]�,��ܛ�,$��_"��7�NH���У��P��-�F���닮��M� ��/�d��A�� #ν���r*��j��Vs���8D$>��r�_�8�yoF?��L���4����,^�I��g���U�����k�h�bz����b����K{+",  c��s���;��hg����Z-��n[L����	��ۘd)�zG�7���|=N�]~G��� �C��IY��]��^+����������NEX��x�|��J�٨R����N�d��KPlᗼ�p����C���H~�7z���������3�~�����gڋ�Ӓ��/�c'89)�pő�F�������4�Ҕ�I	qC���H��|]�ճ���
C�S�7J����Pi"Q�U��NQ�FyzM��ѳ��J���z$���!��~�`3�a�N����C2����`��*ü��F��	�&C��<�������	�����-�-�$b�����9�e��)����F�k/�
�4���u-�Q�aN�I���;ϧTn��-�	�P�݈� �d5�ؿ
p��ly��m�.AV���*�t�s�� x1�{����Foe�:��=p�\���2�PlW����w�b�0t����p�:��������� �o/����M�_�t�Qp�ˁ�@WR���\������\�g4~�o�����s�*�Tԣ��t�,����\�,VJ#������`3,~���S��6�y�>�31ظ}������.'��ܿ���Gs�i�������e�����M��˶WB��?�ݍ���S�tJiI����v\���an�T��Z9��t�O�i����ٷG�b˾��*2{t	�|T�*��M�^�i���J���ySv���%qL�H$1�p��Wi뻒Ų�=�Ep��������������W'&ۖ־U�����Ӵ����sR����Z�K���R�ԉd!n���w]C��5��䷞���2ɋ���O��*��5��M;�g�
�T��k#��Rbek����,;N��K��������΢���}1���nu4IRU �I#�V�WZ*�v���jy&�2-�xkd�,��u���P���U���Æ³ �Cg��qc���Hx��茄s�/���2M�l�4=�qP �rKa5'���	*I p�]xa�F���Zq�ߣ�1�؆u�9��\���9�b�"&�n��˪l�Y�ٖ��_nأ3s\͵i)��11*��iPp(����/���6�^�1�H:�#p����o"G��ccL�gj��W��phFJ �����y])L����?-,j�!m��=���?W$�[\��7j|yR���R��������:6�,	m�W/��ߛH�yT]��>uB����`˷� ҟd��� lwf	���oBO�=�d��Y�(s[�_���)�B�	Oio�:#Q���H�
�8XkҲl�{�Ƌ��h��]Pxɥ[���z<ɾ�˺ ~���'�b� GSq*����D��Q9�W���S�:´���2D>P����Y	��QLJ\���<�dͧ��h��/^���^�f�x�\������&迩=�f����Rҙϊ~�l&�Tm��[��Z=������[��Q����Й��]�/��=�=1��ټ�j��7�m����$�	6�a��i��D�]=^5b�[�#�>5�~�s��:Y�}�l�	5ԣ��>`����%�;W�;v\�2#2�_�x �_�3�Hr~��ȕ	�c|��'�E)O6Ӧ�d�F��G�ZBδ�T�\#�E:�E,�+���1��H��1ӿ�g����U��[��B�x6��g{Z�5w#�����" ���������R�ʾ�1���uwݿ�"Uك ��=m���~�rͨizmw�wKٓ���`rx�6��1��uW����u cfx��"q�:��}LGp��X��r���E�t9g��뽲1���	ũ��)���"ڟ@Y�G���8ua��,S�r�Q��!�Zb������+���l�||� H����#��ߧ������]��5Dݮ0&��F����꼔�j5��@�Y��$1ɚ�<�{�ok� �6:�0#�����[�/��B0��Y�gs>��℘m��sa�]�@��M��|��ො�D�o)�>�*��WWs!ߏ�ܲ�ѽ�p�y��H�Vv�&�W$�I;�_Rd�,h�G7�Q�yφ���{�o5�6��} n�-�|Z^rFA^ā����jK1-�n�5��s>�Yfē������A���-V�& ,���!q�d<1����@�G��	1�ew�9�GN�g�kƜȾ�]��Pצe���SF�[������U�d�zU�7�������n�6JU�o0�S�U�����L2	�qYā���7n���dԨ���5�b.��p%�K�Ju*1�&���W]��<�'���*|z�|��X^r�-���$tbK42����������:88���n�mT��2�(��g�峒��)tq��n�zF���hpp�Qg�UC���ݵ%Z�B[�f���܈���>p= ��`)��5Y����HG"��s��w&��)����Q?3��H�[��F<�ȑR<U-�0�j���~�K���P�N��}\�ti�9P��
�װ_X�����/��ŗ5��%R���X���Y��5�鈝y4F�\m��$?K�T �DQ��j��M���,Gwr��,�x�	N���4k�a�L]�v,�Lk�.������T�{�'��RW+?�ڏ��TH��D� �K�����ۍ���ުZ�s����T�R�����E�~Ըz�\�:�����5���B�q���N61���r���Gw�btt�e$"'I}a��EύK���P�'b�bMK�vӚD�Jr�55n�ʳp'����Zc�I^0ݝl�@}0�����j�8K���
��}-��3��Li�3~@	�����:Rn{l�/���Cu��Z��v+�5�Sp��ܵ:�g�EEv#$Y�yU����@;7~{��V�G�5��������.@[��q��:�e^O
8U�g pA*b�^&�����1����s����Z;FBfdc>2�0��Xq%�? ��y�&���/��n!?���î7�ϘO��&,���`� Ǵ��0��W���������|Io�l�/��2�/l�:ˆ�9�ul�o:,ð���lT��ㆼ�`���aR��"ߎ��|�dd!�-�.#��N�=4�PO��gD�;Af٢S�Se �H��SHo������h+�m|KpC`�2p-r^C�}~C�oN� x�C�p��"������;r��*��^�U���U�e����/���-���" x$�R��5Y��|��� 0�-�I$9����dU^'��a��g'U� ����n��[I���.e���@#Ȑ��A����#x/�y?�L�^�@� ��[�W�"E��'e�w����۪c���7���!F^�VZ$&�ј0Ѫ�yȳ�l]�2J�ި��R#mdW��V�;���'R�e~�D�������J+~v�}�INZ�gIBO�������,��	�8��> hgZ>�ψ�g�ʸU= ����v��a�<�9珄3?W3<����Odӯ�z�XfL1j4,Jk�s�� ��t{*Sn����\�E�v�y`��� eQ���`g��vsCˎ��j84��@gF����:2��Sj�2�h����a�����@������aN<yYM+=�~-��)������$/�VN�L'�	���eJ�wc��/UF:�Z�"�0 +���FV�f;<���0?ſ1.x&��'��>�8�D�ȭ���x����$��f�(�K
�x�.VF���ϥ��W{�*�1.�)n<9�Qpow@P��u��R+�gδp>n�DYmRmc��L3m/ _݈*d��I�T��=谶�`��@���>�l�_<�,�*,����5���B�؞N�%?���J{��Iqp�gzg�"����L$-������F����@�q���h��=CX&8��~��i�O�T��*3����I0��,\qks��w��y��Ja1���\|�P�|f .z��~-.��e���ݥ����i�R�;ԛ(ߎ��oކvM���`��)O�8���z�La<��M��<�������s����/Xȯ�2�	\�	�ު���]a�|PC��hdi(���?�Ϝ Fۂ�9�73B!)����,-	�Id��G��(�O��y[m9-}�
��_�&�X��?/~]���Ɛ���J-�S	-F���c'���r��]��K�?1�*�kgaTB�
+�3��D�N.^-,�N��\db�r�=�uǌ$�l�F�">ؔ�p��'�w�$n��Z�9ԖT�7wmV�B��\��T7x�J���|>D��<f�M|�堟Ǳ�gm�xH;K�49�B>��Iݼ�LC���<=�.+����kӬ��F�q�^�lB�r??�bO�5��U�D���)�G�#�-L����=��������T�'v�Jn~��B=΋C���nQ|�|�M�'����6'P�t��V�����E⊫�?۬a�m����=�;����VEw����= �YOO�� 	Sτ)��K���t3_RH�q5K��9s��5j�lc&��~��_���]���f8nl+���%��O��Z��:S)�ʉ +*��	ՐH	���j漥��YB�Z�\�xa�Q�F8��:��$�����]VU�L>�r(tV�I�;�~��S����XP��A.��JԽ��	���F���wM1�,��Cͦ�7����(xqǳ�8���r��R��z$�W�?��*C�7����Iwog�K}�q�0�3��3ʑ����W�S�����	���l�����fT/�7V�4]3R4���(Aa���.��FWDm���f5E�ۖC�z��٪��	!m^�"�� *�:��
�.�����M�?x�7);^��������2�6�*�;�r�|w�����pO
�@	Y+�U�Ԫr�	VGFG{O�}�DB�s�k��Ii�=��BT�o#��1�Tt�'�p�*jZ��ۭWT�q�+�^�����#}PC�b����ƻ�����4@�'%\5���i]b��`�Cro���)��v��M��6-�����]��c�
��z_\�b�A8.��b$��V���;���ŗ�N���tF#"�����h5�kU����*�|֙
S�癔܋�ޭO\!K׉���[c�A:��U��= \!-/kg�~�F�ED'J
l��q-�=���j�| �"��q��R�]�p"���7���/�T���]��SB�A�g�u?�KQ�E�G�S	&����/������S@�@M�&/����s��;��7X+�~y�nK�KėP�l{�(�q�O�weH����\
����N��})�o�aU��i�h���XѴ��REM��?{u��K�X_����:��i�&�l�]�h�(j�_\��BN�Xd���X>�������őj�\�9U�Σ�/4gZ<�F�Mg�DD'&o[�?�ur�G�x��T�g/�7t�t�4Y9gq����q
���G]n�lst.~;6`?{��ʔ�/S��#�%�
R�����A��re2�H�g�ڽ��.�S.��-D�VU���!R^�"z8�Uר�|����n���%�>M	 �����6baZ����rv�XTM�Q�{��FwmzS����^�35ۥN��L}����U��LοÂ��)�W�����n��'�T�=���ؿV�V[��!��m��b�~~\��Ӂn�(�O�g�{�{��Vb���%��2�༯m�+�6ne����ֳ{��S'���&�I����s��>��'#�x��C�]�Ma�2ޑP��`][�b5�t��A~�'���hW���A��
����w������ >��򩿣/m`W��ap�3ȧ1�)�l!a,��3R�1��pj6�������ڏ�q��=�q�� 	�X�@�> �X��4]���Q�xj��)ϛ34 {��x��N��A~�31� F�/�A�����m�o�m��F�i=dK��s`��K�?h�Ѡ,�*�f���������$��3��Y����;?WX��|�yb]�'{r���� ���	3!F��QI���Z����&�����n<�%�N���:(�'���ne?�Ŝ��z��� �.�u�����CE��χ^�;�$|���dJV��B��e��Z��)`�w��^�O�4df@'�Zd�(�!����²)Y�Ŗ*ԉ&b�&�i�����G�:_����M��,pz�K�s�"K�0����1�,xZ�JC{�4����sRQBi���"ǳ�ڱ0��g�!��E�QW���Z��:B�/��|`�Ɓ#�/qN�T��8��&�L�p5�I�	X:�5M�F4��s>�~b[�qǢ�	L�%���l������\:�J`dO8����d_�[e�d�,1}���W���${�i>��)Ҹ�
���4�d�#nӊ��Ӕ�B^�-��Q�}]��=h��;���jy\{��w�^I^k�V�f"��	��Ǐ�&nZ	�� ����ߙ���V�}��eb~�}�0P�o:�έ,#��(����#ְ#����)�>P�iG��Y�����]7��K�]
zu�H�p��JO}H29���(�U�g��f��/����L���/ޛr��C��6��sHN��Y�'uq�R��G��~�]���RC�_7��*�-u�����>f �aGg7��˗�pdݘ�l,����:����e��+��mk�r�>N�.���;�6�V\�6����#��o�"ǡU|g�v�Dޫ��Jye����G�UE��*��<����*���7R��THi0:�E+�qϣ�:��7 g V�O&ƬO!c%Ԝ���a��Ƶmi�xa�ҟ{l�������nЫL�B'���[��Z�
���l��.M���B�I��y�#_��/g�W_�z�S�e�5]4���%���v�\A��hL8���f���.�g�ʿ�@��}��gܿ0>C6�	0G���{�)^��V*k����C�є��|˶�R�_|���Z��Cz�!vS�eM�Iώ��LV�W����M��>��)U�#^�׵� h<Ѧ��8͘x"[������ł�5+�&�H����c5�1>Θ���B9�W|7�������ٲt\R�p���2pkB�O�pʷ�-|�*X�-*�r�_�:^*��鈿�V���~�@ϝ��c��o0����hO����@��V����h��&t���G�K~2�
g����V8d�Q)LD̄�_��h�����?��������ޛ�_Q	����8ҷ�f���.�RF���bp�!#�O���z�֯1{r��jLx�� ]������
/�&���@M�E���_u����3/hS�����A?��`H,
3aN+s[�G��~�)��^�_�����x-A����6��e�kry��$��c���6DI�?q��-d�@.Cn�=ܘyQ��&%L��A�	71�{�qj/����B��~����}ٳ�W�S ��� ������Qm�3c��_��ڶG��������+3��Nv��9�Ó{�O�u/S���4w\O��?�` B�\
ȝHe��3X #�R�6W�[�ap���{��R�p��3���|t�l�7o�i��Ɛ�(�v��� �շ�����I~g�$𝍁	�ζPG�-��U8���֘�e��`���W/�3�/�}+�ñ`+�{�	�H%�	�2��yw��2��3�X=�aȳ�`>�G�#�\JqLb+v�6(��Ѕ���Lwsez����hO���y���d���I[�Ӊ�,�/զ���3'�a���e�Y��{R0��Xh�������6�"��k�"�r�R��`�qS��g�����U��X[ �k�=�h�[uz���Ĕ�����9:�{+f�y�ga���GTp�.��6��wƕ�ѩ�d|�ήAm7ԧxqZ�e��yq�g4C%!L�~�<V9�CqvsIdL�%8wղ`�	���  #�?e�\���$6`�]��%�|���AuNJ�������OE�,o[�T&�6d���=ߙ��h��.���j�6����3�@˵߃�����\��F�u/|(�1���!���Է�I�7�2��}3���Z�J�؟P�8Vy�ْ����. 7��;P�݋aHIf㟨���@����+�/��2�̔�l������9���3S���?��E?�Y]]��DW��xH���������n����!��ƞ�
�î�dN�Q?���-���Zє�����o�ّ�o����ʖ��µ��Ym�7�qm�*o%vnH~]����:3�WB�V`r����1�X�1[�9�����}^a��LoӢ����_�3��%�+A�����	���x�OE��M������`MU0�M#�#6���|��U#�ǚԐў���[&<.�K9L�i|vr��R�m�{Eة�+ڞ���楠��tD� fj�KP&�V˘sW�L�.(R�e��<��d�T�z_�e�d'u�����|<CV-�{�RDH�2'��":�N�6c������G���r&��^r�qo�M�����[+���v�o�������]����@����a�t.���:�2�sC�Um�C*��u�����	�z������V�e�M��tN�����x�������>���M����N�G�`'��P|HՏ�����}8 ~�Z �Gѷ$v��[���HD[�jZ��-ne�$Z}��fF�i�f	�2��GC��ď���Tl��\m]N�
�Tϰt��
�6�� v<g�O�ȫ�R4���N��Ļ��o��m>���К�@�!�d�Y\Ԁ�U���_�Ab�_X�:r�eU��	���sB��)�9�.C���rc��Sh���l$����n�Zb�껈;���:�;���e�d���s$��Ҥ��3�5
�� ��Z����>f��1 HuIlc�i���iÃ�#R����������%����/j "�qk��&�{i�%���D�[�+��gG[c}�3 ,5.]:�K�Tx��<�����zk]��-c�>t
���e��n;�j�Z�0�5�����Z$1��#�f�sQ��q���ɓ�R��fG�Ii��o�n�����YD��6ճn.39�*�ԇ;�н�}G��H�ƍ��'_����|��PCV���U�%6:�Tq����V��c�$�ߚK�¡����j��y�7�d�DA]��h�@�q7<`�&��Gks���T�f�Y� y%�+���9�!Un4�x4��H����x�q4 @���f^0�2��T�	�oQ����O�ժ�+�	T��zM �>g�VW�Bޛ�X��Ȳ��}A̭�=�|�O�%��
����~�}����FH%S��k����6��o���U<N�����o��:��;aQM����4r�%RA&����Sn�O{�!��*L�5��o�HoB�zށ����x$n|Q`R���`�������,�J�a��	s���;[O6'��srb��H[N�Zv��S�?tƙGK�\��bc�}F�t��g�8��s,�B�`��C:��W���'$�����Q>��/����]��VF<�,3��q�Ʀ�
de!K��sT�p)8���U�1���M��٭�}�.�R@z H���T��
�<i�A|p�̷`\)��Xߊ���!A/�T~�K�֝Š� <����5�ˇd+�k�
�S4�y�}���][��Dr���hE��VEz��{~y�8]������i�s)�^N�h�d��T��*z���pp���S^[�l��\��w�CҢZ^pL���E������s�:��5������Q*��I�PK��:�xҝY�qQ�����\Ҝ�x�7Y���qy�2t}����N6�5۔�w^{�	� cۙB�s�_�I��:�i�鈤r<�O���5��0	O��.�	+����m��
�'���a,� E������G�0�����_Aa�/v�K�R7��v��WHNqCӑ�7%�R��W�__~�ʰ,���Ml�
�G���> ~.ƃ:�),Y�#��Ֆ�0�]�6�/��NQ���=Ǫr!{�1'Р�~R�J�����k��:���ڲ�᧛rr�_�vvל��Gک�\�0�b�jY�7V����+�d��H.�0�v��8d�v�t8uSż�P]ok�	y���;u����k�/\��~��V]���Q�k����:���EnM�-���y�2��$E&?��;�|Wa�h���~Cbf r����aX�Rl2op�r���O��=�b���6r(�����*۱��%9�^�P�b.�f�+�7]mٜ�$�*�د ����X;dØ}�Mv�
�*Q���8,D�yٗ�Ϣ��2Lc4Ci.��4��>���]��0�m�?L� ȓ)��m4�7�5�W@\�����~�F�����x�w�'7B����\��*߫�+m<JU{Je=<.Y����)��+'�3�Ӎ���ɢjә����ξ���W�;X��:9�����̂���Ӈ"F"�*'SGK�x�u$���/���=])^�h�-}�&=�:/�=��\٠��}�� x�o~C.�\r'�n3�8��E|-KV������4_И� %��fy3���Iw��[���(����kHN���P�'&v�Lupb��M�`y�&�)��4�ՃG�? ȴ]��;�ۿ�u�S7���G��~��Q�����8K0[YR�=�S/��}\�9��op��Lߢh/��u��RL�v�J[��� ���v9\88���p�>��t��W�D>�#���Ӧ.�~���T� �}Xek"���d 2xa?��*'���7�8�i�ZWck���슧������l��\�u��X˼z�[���8�eN5=���ߕ�J�F��N�n����S˶�l� �#��U�/��$R<ěy{X��8���w��.gl�Z�QU-�����\�-��ܒE�'c4�#�]_�q�)����$||q�xEL����譋�o����D���V��Z%��0�{� *B\���;�؝�k
��X���憮�=�]�5Ό�~w!c�Ҧ9�q�c����Zn��g��t�O�Pum-���wߖ_���S�i��x 8�vx.3�H{^5n;e�k0O���?��qK�f�z&Z��gk]�
�p��$I�.��ֳ x�cQe�}Q^i��d�r�G�ʘ^㏟�jç�,ݳ��zOف_�	�T(�'6�Y.ӯҨ��l�K>�7zI�P��	����n�3崹�Y��a��#�*���p>R��@'+��<�K�H]��MU����{5�� h�u�t�7>�"`eTR����~5a�~l��Ӥ���{�pL5�T�v������̢2���5ZK��_~I��2w�30_n�ѹZq�[�H�'�Τ�-i4`��`����2T�\��>���՚*�?�.C�8vDs�|O�f x�#/	�͝}���hA�Xd^�a���̝˨�}f�"�f���q˥��ح����9M+�����Vf1�uS�Sv�+����r���jni�����3�V�'��wo�i�q��uk���Fd���C���Q_m!NUm���/������zױߵ���i�`�����Mew�>�,��ܷ��זX�i�`����Bi�JΚ�'�G���r�NN���FO��A�T"����d�CӞ��^5��V
�p���X�@��lH�'�8��;D����l��n�9������~W��Q|%p��H3m=dR� ^^��k_[^��D�k0X��~�ي�Δ)��YW��E/ ˤ�#��u�7���&2��q�G%~-�����X�U�[����j��y+_K0N(�����')OT��fVC��E����
��ww��!j+�����c	� ~4b٠&(8}q����0^���ލ0��� -"1ׇ�4���=�g�ݧ6��[>�Ӑŋ�J�Q�J�h�}G�Ϧ��I��o|l w�\b�.��g�]̤�D���x�]�Up1\��3S��$2�n/�+H�>vM���X�6���.�~'�r�2&+�t;�l@a����b�,��*du���C��������B1~�(�S����
���r����i:�'D�Ke�<��_�Ա(J�.//��_�R�����z��*r�N��{ߋ���Vl�p�־%Z+����J
3��M/�D�L}q��~�<�.F�h��ćd6	��i؜��(�st�,��A�C���|�y��8.�H��(c(��O�`��[�K�*P��Ƕ�?����m­���u`�1F&�/��l��d�{�.[>��� &�OÞ�����c���ayNU�Tc�HΕ����=�㫌*���� '�G�Z|��8�ν��V&�^��_��yzU/��o�|c[>=�`�"x"g)��%�K��_���k\��y� (��Ѡ�L�,�.�ON�'����x^ �w�(p`-�������r��4�UҜ�9��ȵ iL�<�l=������HT�G.��}R3�;Ϻ�<)�Pl�d���� {�=^NU��YS��Ϡa��A��03�"���C���3�v&&Z6�0�{�9�d��t��t�Z�V�G���Vm�]o9C��E:�U(\M����ʨl�?羪lXٿ�|��d�*��|<U�I�K�y�q�B��¡�����d���M�h ��-R��xkw�/1y���e~p�p�H�٨}p�����"���BW���ܽ���Q�
!7xqƞ�.R
�9i+��.��
O*(����Y9���?�BB*�B۬�H���t<q3����5i��"��#���2_Ē?�Qh���8�k�dm�4{����[���N��<o6����&�s5��0�81��߬�w�5��N.���^qg]�Ouct�\�9�X�l��t�\�2��:|�A�#�UCd�>t:��Z5��	�9�u��xD}	�ya�9��h�|���/2��c[�x1�n;��39OBPR<��p��E%3��dO�k��Ϋ�P�䏏}%t��{=�pt�$�15"��:'aEY2w|�? (�SG���P����E��G)�#� ��[wr��n��h�'yX�W�p���ao�vθ����O�[V�q����q�\���H���;�Z�5<Eϟ�
9m�䬛�N-����EJ�r��	��c�7��f�/�~�g�:��r����\p�����/zg�/�[!�q~T���HF ���@����"�R�g~pF�m��-�����8fT"�����>;��_�<���'�H�����vr�+�RI�!>���i`��i/��/�l@O�X^��q��A�^���!�D��1�.V��\En�a%�d�N&-�le�O�|x}����*��UP�����r	2�k����T3�u��X^�j�_��j�,N(��l9�L��[e&�:��ٟc��κ��?_}\���j���8���g2_��oW3�6W���ps����H�x�iD�l����5�+�N��M�{������hm~�Q�Ɠ��#��"stat(8����ڮ���.�ܕ����]"S���G�f��S �#;n_&�1���W7m��ɕ�Ν�I�PSD2�=$Ʀ�C�?��%��(�7B�����M#D�|� ȯ.K^I�_��j�l��Ye $QaOʿ����J}&��ӫ`�*���K} �=��A%G7Wy�χi� =��#��<̠��^k�`�'e���Ne��G�Z�f��IN�z��|�WC��+����7�-ɓ���NG��叼S����tǃ���T��ۺ��SF��������=~��͕�<��QsuU����%�3�q�d���j�g���w�]�mM�$��D�8�P0?�p�ٜ��ĪѼ���i�N"�����2�M���-������j�;����~�ȟ�c� �K����W9�"qK{�Fʲ8tim%ƾ����lQ�J�?:���V�]=Yˬ��p>�lI�/"���[�g���EE�H�U-{î:����͉�� ��d�%5?Uo}�_��r�%�T���*��c��L� .�������~wxR���:�[֘v�)�;%�Z��Dv/&��BZ[ r��6�G�xH=��Ac�O*~�a9reg�3T�OO+�Mqʛ����
��`_6W`�� �8�TN�4R3'��U�Q3���Ot�"�)H#��%4	����u��n���qJ��'�&���K�ru���{����ɒ�0%ي��PA@���rE���ul��'d�� $/�����C�H[�E��<G�>��/n|y��"��T�Y�B�d� ��З�iCr���eB�:�_�ԯ��8l<a�Q*�jU����Yn�68�=���@�*J⅕P��:�}����	Ka�{QX�Ƕҋ�K�9+R����1����uX���9�0�$Y�v����������Z���ڳ!��Ͳ)�*�o p�c����_xP��q ���F��^���C�y����}|�N��{	!Z�����&�5��V�h�[-z]�wB�a��[䫭�X�������9f�����g�D�a�������ٸU�� c�1��F�gU�5��I�V���d�mXɌPCE?4�%�s�K����b��!�� P�<��7)U��H�
�k�mr���D[K��b���h�v�?#Ǝ^ ��֒EvXG#��CY���L��� Hd�ۙZ2�w]�ح���뇰o7�e���c���o� �;/�gH��)��������d�2ѵe�ⷣ�^�B&n.h�,uo��#�g����?ר�~@k�6�z#�lX�nO�C��c��b�+��z �0KGpϜ�Ў�-m[hU���6���rml��^����;�Q��y���'jJ��;z	U��0���H������c�}⿹y���2���`9���&�o�|b����g�T��N^9���5g��o�A,���M�|�)f!U�!���e�Ƣ��G*z�v���p�\b�0^26�9�/ �=�O	��j��P2[S+���6R�H��J�R���Q��"?�y�e3�fb��g?�ݥ��N�Y�^"?zR�d歫�px/��2|��ǧB��˥=;vN�鵑P�{��Z�ЦLt��F�zto�$� t�Sgl��_�q���Ӣx�S� [܌:��y�(�2�\�cQ�.@b��@��H_�n`ԩ�P�`^BU;?wH��5W�N&�s�Ij{<���@o��i��;�<%�| �.ɥ�H��6��kx��_eg	��b����>ע��Pj��z;��a��@����:�qs��"�q�q���h%)��we�)q ~�D���P�(����<�J�6�ь�*��R)�&*3��"��K@~K����ϔ�&��T�4�_3}�$y���|X�2��ӳt�=�>dKt�<���o�%Z\�Pn ��E�CwF�~�(���y ��pLD��3MMN�b��$��s�T�M��1z'��
����d[�됨�?E�����kb���T^Ʉ���:�.ԃ-��wy�oW�}�J��Qى/�/Oƃ��#��$.�����o*g�/�?���4>�Fe�v������*�@���$�z �����|��:,#�A]к%�-�ח�T���r2�2��e4����:}~QjSa#����<O_��BJ�m�PA�
S��[�<4����?�hWvgGZ�qH��2Y1#w�tX^���i��E�;K��iF�̎��?�Q"'8�����
�'�c�l�M(��|��֯b�QJ`|��[���g��M��#�������P�螭��(䢔�A����ŭ<��{� �(�Fͦ�D	LLc�� ^��A�(���3��R˓8e���)���7��lW�'�!�v#�wGCS�n�k���k®��/�MT����6������m8c��#�e��L�����ט��������������Ђ�i?9�K�Q�#X����ߦK&옪��.�#, �����[`�+�E*����ޟZ��a�j噕���'��e���V�a���\O
�����?���8X.���ڢ�
���w�>e%Y�ʅ���M)ۮ�\kqPh��R[	�Z���~�_���cV���'S�[���fiz38mR�DkG~퓑p��+�8.���u�b2���.ѫN�E��cMQ�VE+w�(��4�Fv+�UZ��f�*n_? �'�3�26�Xa�2��4$řA�� �]I�/�K��V�@�ǉ��
�AN���-}.L��Hތ�0��ɴ~4\�������!�������X쓽8������1g5�v� �5ĭ:��.W���%K�6<����/8f�����Nx��ktn��)��l���/h^�WJh}ڈ��=K�/U=.,��o�����BX�Z9�DnWy����Lwl�D�@zoV����{�w|F~D�\l�&	�}z���ҁ�J���ҵ�v�c��t�b!7y�:e{]��F�mJ3�v�@���uu����0�ƪX�D�xWs����)#�ը��sf^�单�%ף����|�to8�#���2�k{3w=��톴ge��y��������bn}���x�O��,��Ly�����YxmRK�n��Z�eӎ�罈��3��Ml��E���[�n�����
6�z6��aq�7��U����@X��~�WI��F�A����iu${����f9Kx��\�����#g�E��z���7���G�r�S=$K��a�sa��[P8�(�'����g>�:��lx4t���>btۥ��Qe�r���0!��Lka�6)�y� ��A.jWm�7�wW��^��G�ל~�Q����2'���v
>*��ރD��i�����6�Xð[��P����p{���-KgvEB����q�Q��M4D�v���.���^��S����˸�����N�9��H�9'�Jf�*k��sg�bY?�H�&�%�\ +��=4�����X��X���U�F�~)1��N���� ���^�c�O��Ry�+qDu���i�Y�^�&���^���)����X(�'�;ƺ~��Z9���n��Џ�1���e�U�����J�f
R��WS8��Ȳ2zʐ�r����}�b���X�铵:z P_��U�R�����o��H���U�V2��#���c�:�!�C,XKG��1ZF4 ^-�L����!����
_�
#��b�~~�*~�o,��=�rSJ�J�N7��g�X%.P�T�E�?u$d���LTv9�;b���e�_+9�_��lO4r��jc֢���x��k��E,^f-�]�[��q�Ĉ�+]'ZI���{&к�� �L5s�>�x���Z�4F���v=���ن�ɿi��gJ�1��{ |�L�sc�4�[�w������EO���,� �,?�O�\�dA5+�Ԛ��%��l�{k�[�T�2�lHc'���J截G`�b��7Fj5�H��Ҭ�Y����HzO��������`���)0�=B��"���A�P7��䕒�5]�9�]�A:��!���rx�K!i��D�f��p��a
�M��[�R(T
���S���-,#ε�;L9~�'d
���e�ޑ���GƧ1���hkv�j�ֲk��@���mlAF��$�Vc�u������4�6{������.�*��)%a�B���Zɍ�櫃0����e�Z\qQ�!j��ਿ���!6x��D��J�ԢgG��^�e,��o���2f�n�c�S$��a-�	�&PUA�9CA��[	w_2����;$�:0w[$r��W�e��Q���u-7�1���AV�3�bD��a`����_	d.j�L�p�[y0�֟v_���� ��Z Y?��hi~�]��^�k��9'���̪�-?c���g$9���zFbKk�Dڜc��F�r�}��<�+,��lXk�R��{.?@H�r�&�q����A/�n5�vu��1���5��<,Q�W���H!��`�6����;Ek��2��3<4p%d�uj�1� ����<E�w��������X�x�!�x5�����' ���J�I�i�n<�]���P���/���f�-���������y7���G�y_�^폾���HU��ʧ�����`7WK�>�I��!-%F���cb�y���Y��5qo�A3�Gw��7磢a����2���<��(��m�_Lt�'���,�h�����Ud�y Q�DS3�t��Ŧ��nWD�ȕg�p�x�O�۾��V���eN� �t�����4�/Bk���˗�(3�9i�gRG�m�T�0,LK+>fR�+�,Ͽ����4F8��c�����z�ﶴ�T���
��}�\��[k�>���z��2f��RPIHH��Q��3~{�Q(��l�0u���׭��"_6����G1aqN��ϡ����{�Z�C_�Q?YYG�O�1��q�xS6�S��%g[����;jz��w�g-"����nX!D�K ��C��iL�?c41`?��wh��������D�-�o��A'��A2%-�N�M��E,\u�S�Dvpܚe��d�τ�0V:vx��>���pؔ����at6��L�L�̾���:sTfKH��ȗ:cQ��k 3�h�>��殮GQPʙ7*�����c��E�s�����������ݎc��*�1 HX9҉�����i�t��Fݼ߁}v�u��U�Y��e���4��=d&d͵�@�������f�crӶ;AbA1�{&�����b�BjtH�ZyZ�!�Ak�k!˩��0r�$b�ڢ�7�mvXmjT�Z&U#�q��I%�I�~n=��z���4M��W�U���h�p:?3�,��۠�������)�zz��4|��v�� �3 f(��lV�I!$|��d+��t5�	r8�y l����L�vt�G��Y�Q0��$*x��LkЭ���2���U�����X3���V��V�"\?�j����J��h7x��s-=b�Oyb�������1(��i�j5���m�:c�S$��,���\[�\����
�D�b�����������%0[�3���:o��3�:��^C���o�C���Mu��U��TΆ�R���^�ȵ8[;�B)�8�V�ӌ�sBfD�L��D�4�ڬ�F�w)���v�H����r���{g���|��ໆ9|���Hs{��̔ġ)��	�^��f�z�꟨���&O�{�81�y�ťC�ձ+�M��=�,
d��{��?�@��s����'XA�&���@B<;S�0��� ;��΅uz<�%$��V��s����A�4���e�J/v�\�V�����>U_�4̉|v�R-d�H
-iu�R_U�����{|��8RR�V_�5erz��g�O�W�c �JeɌ�#�[W��(�4ف�1GTZ]�rE����/~Z�M@>��R-���/�y��/i2�K��j�ˏ����o.�VNx	B���b 1�L!�$�� �q6�^�5OW��}��D���?�X��(	Q��L���Zc����>���h���D������3ŭ�����Q7�7��+JM�8V��e���b��y�hH����F4�	�q>�?5&��d�A���i�_�z������a2��0X�DS�y��6i�)� J�@�� 3ޠ�CHUd���W.ꙤIPE��j�QJ2�����7�?���H�5��oW�@����o�
�	>GXmF<�t�?����E��U	;��;1�M�\����ݓ���t�?֪�hq��x��3�V ��6�S[lF�ب��G��R16>�N��� ���T㎥^}R��߉�Q��Y�4k}ᴣ�!�2���vI�݄��o�m��9�c��<u�UG+Dg9R�XQDBW�qr6 y&#F��e�-���M!d��4�&���X����IQ�������w�:� R�_�o{�KT�o���>$u��"�lՀ��9U�D��ybH��m�yu�?��િ;���_^tp��5}�b3x�ҟ�E��¿��e��? �g<+N�OM��ꇎ4	U��ȧg��\�SR�	 g�O������s5_�ny�T[|��%��T`>�\�Xv��
��"A��ʆ�z��׵C�˨Y��@y��FUY^����}JU�ZDb�x�6k GAB�lpb�`�ug]f��R|��v���	��'Ѐ����v��4�h@*��m�� ���U�줞Շ���zmU�B�9,Z�ޠ˷�������t�h�a�ni/�s�]YJ��&v�P1׌�!� �g�^��>t���K�A��)dB�e� ��>G:u�s��������eWAO�\΍v�R�p����.M �d�%�5�+u`��d>�����x8�R����|���!��ON�
��
áj9��Y$�����UR�d��bԹG�4��;�"؀���-�lɏ���I��Ph)ow���΄��3oW6�yB˼@#;GJY��y-ӇWC���%7�W`��ef�u�m�o�T�������݋�*~C1�0=�q$5k�ف[�6l����VL���<C��<��fA�w��mt����_����U|n��&���������(P�I�;5�F��B�)ۍIx��iw�����ylc�_���OY��
�����O/x������ϴ;'�Nq��E
�M?KR�Tz<1ȧV��f��u����t�����<#.yP���Ч)�w�J�#E���j��Q�İ�کe������\B�q1^QA��$P@�mts�,Jj�_��'����-���R%F��툾�S;��mC�3{q�*�=�U{"0k��&�f�l+��8��#/�����4��K�e	�(ä����a�-ݶFL�b�a�����`~��GBQ!~O6�Yw������@@�Q���I}�8��w+cdG��bt@�H^M��*0��>$ol^�M�PB�|�1�g�s�%�&$�ů��A�����+�wN�m�ɲ�cYl?�#�4��2ŕ�V~zh�@�h�V�}�6e��-�o�Y����X�#P��H��K9�|�"ܞ;� BQ���C�1��dk��[z��8��Cmb��<�.��w��BB�a2,�$O�sP�א/ЧWN����Z�L����3�3�+,s�x\���H�#OH�Q�g�+'A����@s�s��PQ��[�8̑�a*����tA��.KSНͶU�e�	�Y�� 3�*�B������~񞫇���s���#Hwe~s�Ž׊9/Dr%�9q~C����U��iY���P�O�ts����S�&���Rg�s�����y�|��7��)N8�)�Z��I���r�'��b�{�MP��L�s�o�V�Kp5���_;��S����?,|�2��5d=�/�!| 䪟dn�����;����w�UZ��r��5nV~��-�O��q�|S�/��W|fV��sٓ=�����-����/5�Fp��:��#����t�iX`3?�耊�¨nЮ�������"b-���^��b)�R~�{\��N�Q��P+M+�+�Ю�e��_俾 6�k%���O'�+��c���զ��qF�FW�}��Kً��������n����>�;ӳѡxd72�)b�m��t�A�i�H�:,�ˢ�*BI��$�{�&��;D�z_���t�ʌ�yҷ-]�{K?�hR�\]��#�/�F��w�j�S����Br���ሥ�Q�~h ����]�k���=4i6��X���E�+���e>���M	(�����L��nL���'|Q�-x�ͧ�J�J�8"f�ǱK��D2*�,jo�s� �����+Ѝ�3nh5JQ�
�u�h��xjX��6b�� ���u/zf�hE�0��۴����[m�=}��-mx�+ݚ2Wƀ��RˍR~�a����8
��9�	z��L���|�euz�L����`�V����13�ӧ���2��rh�b����Z}���~�� Y��,��d��"������),�1!fĚ��,\���fn�ձ��p��$Ɓ3ǥE�=����1�mr�M���M�qsvV�Ӹ��д��ҰN���L�4#��$4�|x#��R`�
�p=�tU+��Ɲ_^�ITV���X�G�Ʀ�;K{1|���i�t��ƒ�[_�}�d���[mKl�`*@;��	D��@%���1o�����\9�4�d[Aڥ�"�n|Z���K�������w�Xo�K'$ö��ܷ4�$s����yִI���ww�0J��oԜ3�t���B�
�Uo��u����#MK�L� �����x~���O�|̪����Iv������tz8��y NM	�{�� �	t+���x�t�D���P{)��T��xY�	����ʎ����+�p̌�:���TO���j��ﻮ��0��-fœG�� ��LA��T���j�)g�{���P�-Xsm�}k�c�V|��7������#aw�*ۘ�HP���RFj�Tu<�!O��G���\�N������'���o堁;8*��o�ɧ~d�dEѲ����\V�/�5H�H��U���T�%'��~,�/�1ޔ3���X;"s>mh������vl�Η���@|^}Y���%�J����I�ù��{S�X/IPw>+{�E�XK����C5�'P��6��rZO���N�
�.��S�<�����>Y��y��%� [�Jۦ���U�J�!�I��[+)狙�y��� ����)�vQ��>�g�&FZ�\oȯ2��W6L�>��Ȏp�82������X ��ˋ*�Ű��2���xuOy(���y�'kG�+��)���
CXw��;��8������P�wޕz �@ݕ>���%�(�RZy���~-R{��l���U=�iVoB`P��u�0�Ul<Oy ��#�0�%���Z��L�X��|�G�����,�X6%\CIn+P.㵓W:���^�iz��N7�����
���7m�c���c����ǻ��_�:��&=�NF5����oH�������ҡ�wp=S>�7t74�Fν��$����[�W6O}2��XR��U-�v�o� �ո~gVIҤJ쓣���N���K_�9��Ft�L�AO������J<�U(P>7��h��̬N�1P����]n�+��K����X��2���o��m�ٌ�[�j�P=)�[��`����C���1C��G�5`�@T~�GB�r�X^�#d������Ȑ�
���? K�9����a/Xl3K3sM���l�^|r!�:>PYlW��
L�(��H�ؾ�^��&�=�u���
0X�xs�S�RQ�G����%��Up%%,R�p���0�_�O��q��oe�o��c���{DѺ̮3+YkЊ�@��:�����?����-��W��i Az.vDss�t�����P��̐��֎Vq�<�Э����ɀ��<��ݮYF�W���k�#8���y?��B	/�'��!Z_�^��ұ��aع��/&av|���5{�j��WM��6�o]��x��+��Uz�����v�R�C�2�Uw�2�v��1�/-u"����l	�����0�M�4C�1xb|�`_ϩ`����;G�_�`#��#Flb��L��Wm�C�P��vk���L}����j�_���ۑ�����׉9�K-o,���ȸ!�P��<�1֡��s�|���T�����e�2��xi#ݐ��n:������*��(�9���[��Y��;���t����s�
)�\}f�N�]q�.ƌ-p�'?�:��ye�$ӫs�Ӻz%��o�T��wq+��8�f31\)P���t�/���f�g�C���ol,�:6V�m��I�Exxq�p.�q%l�,JZVY̪'�G0/9QA�ŭ"h�|�|�#,��k"��]/��¿2�Y��]�C�z68j��H��<�5� ����d� �ٻ�*������t$�^�| ���i�B݅����4e�簪(�b��h���-4�o��р�3�ڥ�b��
^}�
G�t�v��C¢�VCQ&�:�G���ԿU
��\�0���$�Po���ܒ�����p=B�����:�q�Ğ��+@�G�񄝻��c�,IzJA��I������Qa ]H�lz������&�g�CNQߓ"Ib�@����Tb!��4����v�Kr���C�p5)v&��~�J7��8���f�ϴ�o#�c���,�R���=	��k���ߡ>V���#�$�j�.| ���,���+�> �Ym�G��H�pA�`�g4.n�c��9@��e\���b�Ac�|3O���w��7��[�8�&\��bX�&��|���y3�
�TO��wa!G�P��p��~
�K,ԟgu�;&���C�]�CԽ�r���i�G&�$悵������|B�Ӳf���4��������/���8�赼1�`��V�A\����w;{y���-]Y���X�*N�X�50��mǫn�LY��.��Ȧp��Y�4�j�Ҷ|��V������_1b
�=?������I�C������׿��y!:j	�MN�pH�@�+L�$��  *0�.9;Ԝ�@��d�l7T�r�YG��i��b<����"�Tt)�)C�m���C�Q�E��gj������4R�Ȃ$�ER<�������\��7��'F?F&/�0�2I�wJ������������6jA���8�@�:�؛�~p�Unh���42E���kW�c{�d�D���u9
�[X\��B:��z�!l.�m�!t��8�%��-���+��ȿ�`0�-��v�WY�[og������c���#:�;f(,�DtjY��y+����kI���)�_w���p��p�����+�?̛.�s�K�޴�]�9����������"7��؄��yXa�������u�oN�w ����9R�[�b����+������0�;@��m�/�0�"{V%�DӜ=-� ����uI��m���^�Uʱ6,�QQfqWi	�oNy�?T`'/����'�KtF��wiЯ�Ѯ9o���]�?�>J_�|J\�l�"�f�3���!B�[&ˬq�Ijh/q�N����}W�w'���W�Q7��T�.�;J$i����1H��{��μ(-�������m���p�zx�y�8�n/���L>�)��� ���=æ}�g=�A
��v�M��ޛ��I[W�=���0?'�͈�[%t�[�����Qr������L��;S�q*�F��^A_���-�?Iz��,��^xp�"5BG��q�þ�W�s��xA���4c欧=�W�B�k��$�uL&^�}l�[v�(��={����U)Ar�&�rN�bB�i:�Ȝ�C}�W��XII�jHkW,]t�o�Cc���qK�w;��%�S�zY��><���EK��!�:g�k�:�u�v��o�������t;�S<��M�?`S���\ߧ�Jv�~߃|T�Ϟc}� ����T�&> ?�~�&��PGoj�'˾�T��V��z�¸�J�Q��4qr_��f��[��MǓ7����[�8��K�+]5��ڐR�����MD�]��E~[�Fα S��pl��$�J�����}t��uS��O�H���X5@��M�����
��uc�V�ge����8}����h�Ņ�$�BI���E���N�gϪm����F
o�n��v�03xF��Dׄ|U�{�}<�^�`��i�E�2�%�� _t[���T�b�,]�g�h*�~�'�6E�6}8tT�NL��N��h��*!��,���L�%1|}�Id�	�9�-����mg��F�+̡�Gn
ϴr���9��k4͌�T+�"<<�����#_}ȓ�X�D���o9��N���F��z�QSFD2c.�}����,�릊
82��Δ� �x�VB�c�U^)�`h��$9#����/Z�fx�\D�%t^�րK�J�����`&O�˲>�r��N���_�
�G�1X��*/�4XoMM6���]�`���h�k� �Z�f;XH��1�2]� �('Ko����2^���"PV\^�l�^I�٘43e��M��!A��OԻ�W�O]��\��{glۆQZlR���W�;�ƈ��-c�S�p�':�kc7̰g!��Ή��z@=˳�[54Rn�rV")�>7�����T�6P�o������V�q�
~��mֺs��S �k��?�GV}W6�<��Ej�[#όw^�>�ll��?���[\'��MGY?�x���m%��>���ײ���!�������������C�C�^84�Rnv�~�������=T~�%�ѽ#��)m�8?���(f�E�œ��A$巏��'�ԝ�.+�S+�m�W����cml�FQ�}�4@C}������Y)[����]n� ��oS���t����X�d��^x���=[v�K	M���"����ud7W+���k�c�4Y�
ˍ[�����u+ט�_%��g�3Ud��wF}���_���[՚�-~�W��R}  �r��.�̈����r�E:��n��S�3�S��G��iO!��{��[�� S�xu��J�c]�w;�H��Ϛ�Z���>���,uyND1#dɰ��w�ll���s5��T���q����ћ�7T)�Xhb��r�U��jq�@��z��Of��q��ܿ�I�HK��������hSTB�g���j�F�(^�%�`z���!QDI��8�oc�^I���Ƭ��o���?�*��He�`�r�AÅsp�3�2M�D�"���;0I�rE	��	Vѩi@�3e{��Dݲ�N��z�� ˧�=�=�kP�WYU����1l��!�01���PBPM���Ȍ�ԂN��vi���� Ǔ�o���_���݄L�5��T���׬�au;�L4u�����*/IU ����ǡ���c�**Yu%l�;T���Wv�f�[|i.ќ҈wo%���o<T��hƀ�?;��Z0,b�� �j2��T"Pd�3��'�ܭ7w�c$J�}ŭO���J0��N`��|j����J-"��r�C�.ѣ��}������
�8�=��%�p% \O�����u�X������rj���݊~��,�L��z�Ox��O�c�z�i�Qy�s�S�]���d�T0�� �=߅��.�� ��$�
Q����:E��O�\����=�S���P=3;CŊ��=��kg�>����[q�BR����l�'o��R95���_��/}�8����e��v?CJ�V�����>�Y�wv,?�Yr���L��WK�}��e�T��d��f�ޕ�Y
/.�{b�B��.�����|e�3ߔ����y�
�$e��z���y���ı�&X3��b,:]��_3���WūG�iy��O/&�%^ݠ���||��@GsɆ��R����m}�z�1[�"�����f�6�N��ȓ�ؕ�Wx�I_��e�`�W���`�'�.�P;���C�N��)���1�an���09��%�y ��a����(�C\xH�1�@���Z�.�1��M��\�ے�Ģ �T�S/.*#�dg"W��`sE-�*�Y�z�:H�E*},���	��_�|�V�j�x����;�����BkRbI0
���)[{�Fw^�Hy�շ�m�>��}��zlH���цU�'w�15�\>[��-�����P�b�ZW��J��`IZvp�:��Ew����*J���G8����> �j����dY���5�4ݟ�L"�!�gG�ula��-GR���Ld��7*��ɇ�����/hxK��=-�T���֊�!*��OD���#�A,���#nMU�ƫj W���M���z��>:��GV?�W1�U���*Q2�L�:[{��50���<܇��1��m5�&1V�e{6Q���`�����`J������gu���r;	I�H�Ƚ3sqsȄ[-_�1�'����y�)ix�I�����Ϊ�JD�09W Ȏ]fgq/���,�\�����?�����d;��W�g��.&x�TqqD�^�#/j�HY��'4⟦GsU��/��PB ,��'r�'/8VAt�*�k��H�V8�r�S(0c��@L��Z6�t1��Qe��
��@8�ܿ���8/D	�r���+)��L G�����B�M�a���� ��{���x9��C�+C3���y��Wfvdq��w�:�O&j�liV��4�06������}���rRL��1��42_�S�șߧ]OkQ�zW� B"�f����;�n�.;�Y�D��oK�����l�R6��%�:C��}��i'��SK�"�-��xq�$���<#yեgG�I���ӻ��Ys�[s0p�5�ːb7��~JZ赕�T`/yS�F).�̚����|��f�/%������hE$��'��{���Չ�鼴�,�H!-�l���$��6~���t�]�d@���^���_��1�a �\eAlG39MY��6�Y��Y���[��^;Z��Qʤc��4i�ѵ���>�5C}]��W�~��"��]�s!%���n����n�3IA���\�B��$���'�k`+���q�ͧ�5o�>d`O��T���r�&���0�`潪s�ϐHV���l�~���tE�= ʡV��:]J	�?�0I�%`��s�o��R�>�8��������8Rj(�/;���D�RNt:�Q:��r��1�z�AJr6ފ���ǚ�Й�r���i�n�A�����TڠսC
�_[y�$%ėfâ�E���a�b��"�5]]���g�ƙ9T�]��΅�P�١��ĺ�(������0��L!9���!�>�N��|�U�i3�L�UO?����=������#�26[�[�̪�D�8�tTZ��[��.��ٲ����8x����ij�D��	��۞-(��Dd���l�&�����>W$���5NG�2��b�afc�u.�oH�
*W�	5�`�<�s
�tH�{Ll�+���'s�����Ss����Q��@� ������z��M,��_��Y3�	���B�6�_��	7�!���]��ʑ�Q-fG��.� tg��F�[���`e�LK�胎)S k� p�|���.m���@k9u�h��x�����iGst�e�F���H��� M�Ţۿ�Kܳ�B�Qn�S�z�=�m]5����3<��ն.v�~��HDw\��%�i�P�*������w�
����YU�0�>Q2����=������iX�x��D�`��+P8����q[I���!�ԴG���4�P(+y5\�B��fO�5m����BK ��R���%�hV��Wc�����+�i��d��t��*��+����cү���ʄ�.����>�׉F6��ɒٺf�8�04�`�;?t�d�<5=��"�v!neQ8�ry�~���V��:���Ub/jY���:��hޜ�����3�J�Y���AI�[��րm$�H8<��So��7J]sT-�id������ӌ�5�`���㇮��X��')�vc�����>BY�M����W��\��a"��ǡ��͹I�����F��kNu�ڤ�p����`*�P�<���A�}��IØ��}P�����$��^��'�c�iM ��hS�����9�7�"��x'E�����yl*�t�x\�׻+9M�q~1//u?sI����E�<rsR/�A�uh��K���p =�d������^�;G��MU g7�F����W;N%�W�Hr��3����Q�-'$=�%�
�w��	~�b�bmK����g��nq&�d��]9=2�@�fׇB)�#����w{[f%D����g���>>�Io3�#:�
�F6|g�<�����j�(�l��TM�=���Nb&i�HP�g��{��H�Y�RA�S����&�=4�f���y7$#��٭�h��$�|2��i�m�咇�8�����ѱ��(4$;��љ|�/�ݪX�PF)��׵a��wqɳXlTf��	�O�+?�l��Ã���mۂ ��E�)S��dN69�ح+��_��BB�o�5!���d5�x�<b<l_"C����_�;5C�.�#ξVL��NM8���F�p�ڢ��q�p��r.��|��zC�}|�ۿ���;�|I-��I�ߐ��W�Oa���B��D�|���wْ���w�t��C1q<1�m�0r�8��	Y���b���0�ᾉ���5~�n�ye��L��$^@���?2��F�B���X����+�G�rC�'��0��>������*���mI���m�m۳��f
��qS���}O��N?��h���z�VۓF��-��^�}=q$��)��]U��e�S���>�W��s�u6#�D��D�3��g2v�}O�q��pBD����y�g�[ʌ�b���2:}(,����W���j	~�а݋C��o���!����(�`�M�q�ԬvQ��X4v�bVx XB~N�S+'lX��#|6]�k�'P���,���)�v
�q�D�������FW�@�bG�cf��;��|á�>���ݝN�[՗����� ������B.R��_���1<�:iX�q�aP��>jGol,Q�=�0NV���!�^�>������)�?Q��HCл���]���B*��?!(�d��k�;��e��wm�b�#���5R���R���Ԍ��غÉB�+����G��;H&>"����{�B�h<{nN���.2rx��
����� �]o��$~�O��C{&��\�pB����=��pha��{l���gHF�3��&���.���š��z���&:�qU��@��h���D�А�e}�7o؇rI�v������CdE8�k�x.w�]�gdEާ���v�'�7eh�.�����[�Y�}t���SFR,}�G�K��)K#z�u�X���|ޤN�G�Wv��4�����	.���'@p����6���@��!xdx������jﵫ�%���v{�G�ԏ��Z�\�W��g��QHHC�t>Q4b+\��^�J0��}ɎAF��/S����؍�J�I�^���ht���)O��t�\-�RK	^9��G=v�$ˌᄚ��YJSksu	nN���	[	[x&��Y��O�4-��U��j�c��Ab�;M}�"/6���qE�/�b�N{`��c	��k��4f��)�$�oml9:wEWT���We��:[�k�0�� � 0ѽ/��* U��V&��e�����`M}V�MjN�8���J5���$�Hw�qG��<��R�'*3bZ}S�s��i��(*	��.�]M��0d�Iy@+O��Q�J�H��͹d�;���$���6�?�����q_�ٝ�"ȼN��T�x��ܪ���:pN������T[
֪/h���/ s}=�/�^�Ii/^ۺ���Q�����g�U�IUx� ��K9����멦}i����?*�;v�G7K�W��9���v�Dd���#�H���Wt�T�z
��v�!p!���ܑ[M�Nd �z�9w�M}��KLV��R'c��a�ʣ���A܏�x���� u�٧0q��z�gU\����aL����>��BR_�*'��?��H�׵��=��^[���b��gIӜCʦg�[2�s�g�Vq��U�	e-4^��Z��{ǈA���S'��Y�$EN��� 0ަ�a������R~�Z�c��ۨ.�V��qM3�P��*&�j^�P���
H����P�Z�1��SL�"C��bܔW�ʷ�/�$���N���TO�m��2w�|��z���Pu\�%�Yuv����^!�v��CMV��|Ar�+��;�uj)�=0�7���~�>b�p�T>��|��I<O�ܕV\�Xü��w���Ah���_pf���E�I���L��Y�X��S���^�J���.��z ����/����"���R��K!SC�_�?�W��JU��}!U-@���Rt�;����=ۺ������s��p�ڲ� c�7	�L�ΛWG�rwx��/���}�I�$�����P�W"�hc8���0��Nw�`7��;�j�܎���'qDF~��dmL���	��\c��U%S=:���v�拓�\�;�T*��6 3�Cٹ��VR�ͯ���EC����"Xk�q]��Y������ ����[�!U��EI�Sd�-"z`�f���'�My�.����_a�s>�n<�tzF�̅S���$�U�&��l��u;�$*^�5n_�*�t�\�+3���%��t+Z����Y�9iEQ�3ȕ�_@+�;�����!��Nm"�?�(i{λ�.IC��=V�S�5��W{]�p458i���
�I��%Z��_D3*hbe$vM����
�MxߞTC��E%_Ug�F�5��39}MS �ʳ\��F�྾���R�&����0�/ݜ�ޜ_���!g�_�%U��@��C��!�B����'-���w����_zrDY�B�������t�:h�����\�k��?#F��0D5�D��As�?i	ruw�s>'̛�m��7(0�Z�~�iSɻ�\ôOS->�n�p�5T/m,L�o���x8�g�P�ɧJ[�a��K���`���9tl��6��D�W���e8P�GB�-�t��Q0_~�\�(嘶Q�M��=IK�D���Z[����n܏ț�V?��6o^�U��>Q8��m���K=�잞g��B���H:�b��HB��U>���b��V~��#��w���� �	���t����Q^�B�}v�>Eh�1�/"̢=�a���z-E;��[ec٨��}� {3#Ǝoļ��NrU�K�|�o2��*x�{�A��#$}]�N���N�dI�[�9n^�0^�.�>u����=����+��>�H���ў�L�q<^�Ýz��A�S[&�m�>�u����e`���o�a��o��#0L&�I1���%�u/���y�J~��n�q����LP/H !WI�H�B�{�o�#����n�k����w�%$q�%��� 4@ʞm+����\�Ej&�Uk�a7� }�xz�c/{}7&_S�V�^�q��!S����2��u-J0���=��^?ߋU��j�YT�U��H�Y>�خ/��8��sǪ���3#��_�g㓚R���R�U�P�����7�𚡮��zY��Ɠ�y��\�u��Z}�z�5T�ZZ���ոɿK^�hz-� ;iU1j��t��Qؙ�'Vs� ����D�>+_�~t��P8�V���+ �]
�8HwyX�e딟TGu��D8;C1S��!K�
VeE�Y�f�� �p�I�1�	�ijfC.�ů����&"�z���9�eM��b;'�Z�V��H�qG�$���(Rrp9"*�*�#�ƪ3�%�Z����<��=f?e�6�d0���='�5���&_ߞ �*�[�C�l�\ԓ�&ܵ�;�.RA�Q��>��ki���?��P1𭓻����Ö�(�Z^�����J�s�vRo�c��Σ�9R�<�ꎲH�(�c�$�����p��p"z���E�^�����G*�p f�+4����՟#� ���o�����4\���+�6#��3�(�� &�� m9E�:	Y+BD[_��N��#b�L�:%M~m��@s���7Y{��C�� $��+�5L���xo�0���(:�����z�"���+@@��܆7�^)��Nyz��r�j�� k9�Z-ev�?��f�[�O��IR�W%B�Z�8QҞ����I�\S�ĕ�S1B��+��nD��$��z#l�M$�	��ޝ���o<��q�b��/9�-�^�'���ժ�b�~;z�m��[s��(�a�8�?����� '�u���t.-��<�n�>�"GZ���͵�xC5�]��{�p۳���%P��a.��_>|��pVR�T`��s2���Z~��Yz6o�_�wt�b���b�F?S��"Y��s]��ːJQ2�r܍��9��[_Gs�dX4���x��-���K�7��7��I><��c+1�x���g���3����Kڒ�ȕ�(�8a;��}5�����j=,��j
�����=�eAP^04p�jԍxe.�y9:k��/�9�=�\�F�V�s!2��������*��Mo��CU�p�B栒�	�"��7[!���t��oƏV-k;-�w��j�`�����g�N<�a��鍣�3�Z�ٞի�;��Nw��p�r��@PN ��5�چ���z]u6\=}�@���>ȼ��0�c�ћ�g��U�kw-�� ����l�fDó�����߹p4/ue� a/X���؎|tE�w�.i��U�n>�N���$v�w��{pe���6��ao���1���*�T�[.�?�<.&<)}��1,�	�˘��iAx���>Q�pfJ�.��o�>��pO8w��Q�j%KB�n�k���{^1r[�^��!a�Y%��T�E��q�W	�ܩl2�z��>fI�3��x R�)Q L��dKO���&��/�|�û̇`�ǿ��無���e���Fq����y�8�*��Yf��-�9�q��⊢���,+�Q}\��B��D	wg���̨�����zb&~Y4�Z�g�=x�%I�:��k)�,��L�_�#e�8\]ɖ�@Ӟ��5�p��j�"��Q������1�Q�Z
̆a�bv�(�{��}�N�]*j��:��9j�;|/U�B��P1��[jC޸������@�4p�m�"���)0��&i��s����O��b*�����Fs����<��Q� �t�T��Q��y�'���p�y`w��<Щ=Bi1��=����L����^�x���K�6A���,���6@�1N���:�`���f�n���ܑP�C�n!�Ob��F \𡿋�5[�r����~���ƭ)is�绿ӖgFa�������9~�ʒ���c�w:�Zjv{�Q�-U��.&�K΁1��Eɇ3�� ��֕�}�&�Bm��qʚ��l�*�(����
g\|��3�L�qݰ:�r�5�[�Y�K��� ���1�������v�z�i-̿Ǜc '����|b�<������F��k��5竨�U��~O�l�)C��*��o�	�#4������\Obq��w4�V-����qP�C���F�K��!�O��J�� ToG�dR3SB�Q^xp� �3u7EIA	U�����p�WTݛ5��M�;ˠԈ��՜7�|�&=D�<��oO8xB*k���m����8|.�;��}����}"߲���'9�NJtN�pǺ_b�����T'�r�B�?�Ժg� l�YP|r	��`��	;��P��񇭕5_�Z�ؓ��Էo;��6�F1�G��|S;�[��5_%U\�	?�f+~z�q�/��5�缭&r�
 ���q�>0yu���o8�A�\������PH��͋��7�� _�z8/��wj��6IJ���m�P�wM�R ^S��MXq�Tq���&:R�����#��u�f�E�L��������˦#��o�;([��@������`�aF.ixa�ϝ�OW�D��� �٦V���__�����{���p�Aɷ|���6mpG}.����n�g�N���&�4�����,�[ٛ�;�цnT�NLOCF�!M��0��{j$Ȉvꑍ4��-���;|������f��"�ii{���~I��ǫ�U��J��et��+����8�P��}˖� �B;��֭�
�,�_i�ܾ��~X;�7��$`Y�z�p5�+n_�1�����8����zղM~������&�J��F����G�Lb��}]�s�}r*L�>rw�[��_�;q��e�θ�Ұ��K,�~�/�f4�@<�eW^լr��G!D,.��"CѶ�{K!���~C��3��\� ԰�u-��9dg$C�9���x|V�P��ؠ��G٥L���]�ݛ(���k@���j�`��"�y�%�A�7��V��+k`�W@%��s�)uW����K��� ��7���
{���S�&����풁2&���l�N�Eğ�\�~x@�Hs�����nW���[>>���]���-��^��_[�`�������Eգą����*a~����Nj�[XQ��M�|�Lؠ@�n��Xv��
t�&f�9�<���� Kd�<�+�@�K �"�C���6t��� ���'�z���rU����±c�ǟ��)�
�$�����������)C<��M�˞"ǵ%�}�DA��ݔ�5 �Z�NJ���j> �'B|ǈSr�E�P��t
�7�)U�8�����ڙ���u�@t����R�6@�A�ޛ�}�`�|;K|DL�G`�gVÓ�Z�q�L��ȥN	9a_:ɸViJq�Y�N��)���6[jE#�V����a���\q�9�??�@�B��a���ҍ{�3iR�`J��c[ʮ��v���n�x^��2��nLmFQ���#�G������n�0�� �E_�?��n��o��Z#�������t&.�D��o�vL���$�� ������^`��@����8�[��qs���D#�Wг�KMb�+���L)�ԁ�ŷ��h��<n
��[%w��B1)H�Dޮ���Uoވ����g�&.�RY���ij$޿,!�E˖n_�o���p!��s���,�E�o�i��h~�%�nر�oEoM®�Q��d3�m�+ V�	*_
�
B�m�x_��"Zk<����+�F3}Ġ��q�n�V�SK�S����u�hT]�� �k�x�<���;
��-љ��P�?�>?��M���K��.��q7m�s������e:ݟQrYi%�Mj���+��7�uE�c\�o*86e0򘲝�Ҹ�E�6����	H;�6�
/��_���#t��K&�,=+51_�Θ����M�A��+��Pu�6�&8�U��S��o1%%)�\ ҶN�E�lOw+g�����1Ǎ��l����^��p	��N5�p�N�U��i��CnJY{��a>
צ����	�D&I��HS Ϫ>���~�(ׇ�A�-�ӯ��`�C8v�����FB��Č�߅���ވ�x?�L��Śl���,:8$,=mD�5��[J[�ߟm�q��j����eDWٌiƐP��)O7�g�#<xm�������Q(P�Y��v �k�a�� IjP�;[4�_%X>���g��K���>ڸ�)��*hb_
e4Ce�>��SD�����t`���S?���-
�S��x��x$Q{�4���F���(��E�w�5xL
�� ��~���f�.�JJ�^Ke��QA_O�r����[jv�������AӆHw��W��KB����B�c���E����a���5ڈ'j{����S�B���]��G4W,��"e�"<u�hp�Kj�_��IKY/�T��EHq��D"
�FqQ\\��J�V�PwQ6�t;F���D�V�����=��v!��7Q�`���;�U������9˞"����/x��P3���O$5�������)y����!��tV�e/���y�eU_hOG]�DlS���k��AjكW@��q��f,חuz'�Oc�P�76!��U��B\i ~v���!����N׽ܟ[�f�)+���"��H3*�l�&�P���O��l��b
AQI��!r���'=۩S���ę��}�w8&T6�{�~�����/%�A���Yɠ�����\�j�������B�A�����S���}J���S�&<�⢦?T��Q���K5���.~'̪i6�{�w��F-�KH3��$�|�fR<17|AQ��NS�+�[-"�aeC�-9�ٲۃE���'�%G���k�}�.�3Om�]�1�����5)J+s~"�#hi��MU����g�B�1o%�����	�6������E3+S��HH4&HƯ��)��.�ހ8ȊM��Q�h���=�[bs���_���5�8`������g���1}��F��*����l�:�Ԩ�5���%o ��R���&�������]g��/e�1*��X }�%>�ѻ"`�EݽZ�刈d������	���s�L~Κ��˛�[�m�:5�5�^�];�g^e�O#k>�N�B�I;��(F�>�SCR�Ќ:���c�eL���
OK��Z[Y{��4�G�,3a	������A��]�������#�����ʊ&|p&�U�<+�j����*��y��y5 ��(%��R&|��C������_YO�N�8�s@���I&y�$��җ���D�J��$����P/�(��z��������A�:�T� �;�L�xp�㐿u
����x�<�~�s#���� >pqT�3����x��`t@UW���
hW�U�uǟ*nK�S ��l]]U��/�3 )�Q�t|ؽ�� ;�l�h�������{8���y��g�ح�%�	��7xy2�(Mn�����V�Sp,(MRG��P�[N_Ʒ!���8��������&���+�h��$��0C�����UKԫ�����6���F������@[.�U���S;�9"�����+r��~��M�Z���5��Ѭ�qN307��e�Q%�n�����''|i�1���=���b\>i
�!ӟ��뒏�_	i7�l�8����-u����E���L߆R.�����D��"k�֯��
i��`��aCZp���|" ���N51N��R�tM��ǅ��<�}�K��uY�v㊀�h�Ó���O76-�_��U��?�>��u(B��u|Fab�Sl��90�"��Ċ�}�9���X��7	�_��ө.�,�'��>5�`��w�@a����M�.1co���V���P�3<����p�0��ޗӵ��wE����8L�������ǭّ���e�s���7�l,���8��q���8�>�垅���i�L��8�k�Cw����3��^ovp�p�X�p3ݩ�'/�ʴk����H���qE)S?���;�C#5|B�v�{�m�aR֦�f8ꣶA���K�@dd����UM�ͪ��W0�-�f��}��h�@c�t�eج^�
�G-\���"�ꋎ���r�'�{�|_��t6�_;��-�}`�]�����U'�`]m��d�Ċ& 6���#�M�@ʙ�qv v�����O!ꊉ<*��
!�d��1� O�H*e�����
Yζ��;��%	4��b�RK�'�N>mHl��8{����vQI��^qR��6}K��}�EJ��{%r�O�{n���2|K�{
�{�@��;�<�ꆎ����u)��%!YpP� -@�x�٘�Y7}Xu���?#�6��0�D,��{_ʝ��c�©�/w�V�Y?K�jZ�#;���*n�� פ�Kw_MTH��]�$i�Cm���̮$�cpV_B-���,F�#q�(���Qv�Z�Ь"��w5:��P�Y5�6��O��P�67�s:�����4�R`�?�>�YI������@B���L�4�ZztK��AN�8�%k�J�ޕX��z#�e�φI���`=�]�����D"��b�����q'ݢhc��{�j�(��uHpD��o �����F��	9��;��+ �ؕ9T��������Y�ʫH+9[?��J�����ڔ���	Č-����ܾ��0T�f��hͩ8)�t~F��nI�D���P�0@����V�*����(ewj`��Z!v��q|���M��A8@F����C�G;�K>�$'��F������7��S��OC�9x^ ^ꌒ�i��_�g6��?|��e*K���?A���#s���L%	M�YGO]A�|\	�������͉�mf?N`�~k`;0ȳ,zt{��;���"^M� Kx?hufʞ�<J�_�1�Mةo�����_�c�|�k����Q��&��c��V�K樘�8{����&?wq�hD���M56j���vf�Lx���x="m Hm��)Ф�M>��wqى��8s�-���](T�\�5��S`�C!u��BC8x^�����b�5��w��U� ���Gw����{D<����Z߉�d_�ܳPF���B���pO�P��x7�e��o3�n
y8n	�J!H6ޟ����� �,�pg��/�:�ŗ���2R���2��l��E,��o�$�J�&���?��73�g���*�h��5�"�I�z��&��N)�}����a�*�Ul���(ʁ�IբC�{H,�k�.�!���)ô�B��LRM����4c�,%�F��;�|�;ZiF��|�%��P�ȣ'O���ߓ�E�����ѩ5j���S�e�������	OW�i�@���bL��>�FK�S[��:�;?+s�V���B�_���+�%��I����Ŵ����'DLe��ӣ`=l��acT���}��o����>~�G-��A���jv.'�5^N�G/<�l��u/น� ���
xw��4����`�[}��I�n��GFՐB�sNs~�?�� ����A�{�&���(�/v���d4��בG��!�j�r0�V+�h��U�����D�����>�?�g n�;}��"?�b��\�<��V���;ȿ77p籟�X��_������\-�/O�&���{����,��� md��g��%���\������BÄ��
e��'��ۯ�~�jW�#�Հ]S�Xl�m�jFJ��p�����1��>�8>�C�1��q�my}o}jp��cZj����ި��F3�t���+E3�h������׼£)0,=«��B����M�(�|�GUI��\x�z's#(W����P�Lh�R���^}Z�5<x��j�X��$]��D'�G��{�ц��p_�v�C���#=����
41e4jN4n�#��K����y�����Y�� M���_]�@��-b�ÊF(�k�d��=�x�ٰs��I�̈́����Y8���iE���*ζ���u�M��뤉nxɹ�>��1���oD5��07F2G2��O�o�q��p���1�
��%}ʽ���}tkna�, �ſ	�)���g�Ld:�=s�R�͍�٢����������.�GlD�
z֘�G��%�sU�^	(#�?\�I�b_�V
���B ٸ��A�|X���K>��]6��k�� �ʠ�����l+�R�_�G����Ù".�4� v��	j<�����'�'�P8�;�#,�-�y�.��N���9�NC����j�D&�D�p����&������ػ|�{���B.6=1)SPⱁ?�����9�W�:X�>"L7�v�%��?FTjX�ݽ4=�g��8֬׶o�36͹��c�,��^m��mѤ�g��fU��̒�.��"fsp�nZ�up`�k��5�ZF����flb���BgUg�nG��5��<u�Oz5��nz}�_���b���)�Q��LRY�B���@G[}�)9�ԧ9�h\(��":�&?�4���/�ǈ<O�y�n�9R����������DЩx;���>���E5ޮ3Fg���#������'����*�ۥ�:����Ҹ�!�"8��HJ
 �~e�J�<7.��WXZ�Ү����r��ٜ�#N�/#R�f'�Hbi�j��V������)��Db����[�	(�;�+���wT"�(��Ԅ�K�Ec��}�@��w��km�� ��x�QE)�\�h���2��Ё�It���$k�y7�����=qF�b��7&�&��������8�>�p�K��ir�Z?DC�`���'ߑО��2ѱ��p����'�5����c䯛h�J�R5$�\g��Kw�Zy`,�,W�H�R^��t |"�,�}��j1������3��_r�4�qb���b�|��z����|���4�}�7��������_N��4Ɨ�N���0WU\�;�����O���GAN���0�.��G2�c_�+�L\�����	�#�L�L�y���t��R\@��K�0�r�;q�����(q�ԋ:۩uS�_읕��|����	5����RnU��?�+��e|#����8�o�+ ���7/[8܇��dk��Tv�q���sg��){-gQ9}
�v�	b��9)iQe|o��A�1���Jx���#��w��~��6��j��rw��Y}�6>y>|��o���]S-E�AP�d	�U�.Ż;!(Φ/�Έ���ó��
�92C��uorGQ$v*@�BBi���(�;S�DM�A�
�@/S;���p}�7��P��R]]�Sv�?�4[k���ǡ�/B��W��O�M=K�#/<�a�S#ڴ��V��
�4��ԴŎ��H/q�3���^�+L܇ �͓'�VQ����_�ռZ	-E�?6��^Y�X�x�O�����cKa� ��,j�la��KSj:\���s~ǯ� WA{N�a?��q.:,	������t�:適�Ca�ߎB���!�XԺ�a9p���a������,.��w�@ ���i����J����;�� ��^�Fʝ�Bte��2�`�ھ�n�r7�IT߮�֌����~7WdV4}�d�
��X2ȹ��U0�1Y��
*�פ�s{3:�P��֊�;��9�j?'pA�����G��ͬ�n���\�������N��ْ��a�/E�c�å��X�
R�9�ie�-N���s�Q�}� �B�&*z�a�_��l�h�BE��*����( zܶwӴa�(Ќ�(;����;Br)�+�����q�*�ϟ��+a�w�
�O�����Klf���>Q^�<ޣ�1b��+�Y���Sn��Lb�!����o��W�G9��P��XrlnN�k�z�;^��Y���5�&,{J���uܾ>~���*y���'��I��5�YR��	�?i���������Z�?�ہ���e��ɂ?Hl��oT��ҍ���j*�31���
�P�{���а2B����zq����`����ONg]�(�,��TV��4��
�Ό���@���Ҭ8��(rڏ'm���纫l�����3i�~7�0�������j�B��dI����Z��,j��v���[=����7qZT:��6_�:<N��[��A�<+�>�h!S��T���S��vLD���3���S'��޼ ��6�3iF�V���×M�/~�.����T�DP%��J�סWo')O�E�y Yծ�b���Y���t��$�Y�����)`���I��]J�Ki-wwh����u~g��^����;Ů�X�<�����f��:���K���䦞�h_�X��$=|�2�rƊMksK5RS]Q�-/�*�=�Ցv=lep��ҙ���5�6��O���S��Y69�W���9��6�J����,��{��"U8���J�J�;�� ��W@��u�j��$����)d�^��tq|@���#c�|�qIio�y=��֎F!᧴��h�
D{��D�N�3���3*8��і/��\�� k�����k]�9<��V���yt��5����I�<�2;�m=�K�+�C�Oʙ�Rݤ��?�O6@�j-���"��z,�o%%}.����94�=u�S:��������A��&�s$+I=6D�A�.��F�W@Z�(VA�}O@�������9�O�n�<Y����d�R�)�H"���y�Ѯ0Դ"��_�UW}��ɻ��kh_��U��$k���I�R��U_�Y%�-�d{5�uf?J��Y!��iG1�*D�x7�fK�#,�}���ɯ1ZC�0����|E���bz�('Mͺ��;�$�85�A-�03Ύ4�=W��]���4_�r}<�y5�`�϶�dM���3�T�W;$�x�G�� �aq����ՠ�����n_��ҵ�Ƶ�vʊ�:�%aUN�i�}�1��Y�|�RL��ie�ݯ^V�ߪ�qsI�/���x�-�c$aP��s��2S�rn�u�S���ڑD.T9���2�Rq���)��}�ZԮ/�9�h;(]ŷѰ\ɰ��\~2Ĉ�b�k���K�y��a�_�ǫT������8�͂'��P�%�E���![9S�%��Q�F;��Y��|097�Y��L����*o�j9?�MK��~gN���EM)J�F7�#tO�B�<_�i+���0�x'����x�b�j绥.������Q{恙������ZU���f��f`=5:���3N�̚��W�Y�U�����WZ4:���-�]g��i�"V��Cz>�F��y�>zOb/��!���(�p)��;"��P?U#���M����֧5�Su�m<`��L2���V��m2][m���n�6���Q�|V���Уr��!�o�C�Y��x1
V�(�'@�����] ~�k�L3�j���t ��ۿ� ���ܷ�U*h.l��W��w��r�s����/V�v]\n|dem�Z$/1���֧��&o⃑!��%�ݫ9�1��a�_?w��ҹ։�.�Ye�4$}tRJ�|p��\�Z�L���79y���90���UHK��mI�[�9N�<�=<���s��yv,�ҝ,J�/H	���R2;�	��v���K� :���*�t(ٛK:���%�.Ջ	�r�C���&$�x"4S^2j6�sl�����T�b������f����<��D������X�7���z[�bc�t�b����NDV�e�u�!��t^��k���[$��ޣ2ax��v�ԙ�|��!�gRKR��c2ъG�'x��b�O�ߟ	���5��L\s4S���1n����P�w$�Pr����8f���-��l��1�aJ-��J���h�<E�n���V�{Rō̉3Q�"ڮ����G��7~����
I�N�������4F��&F�l�������w$>��Ydf��l��ֲ5��x,]�ngNY_gg<��[qP_��.|���b��4p3N��qܰy��m���|�kDj�/����$T�BϢ�>�CC���}o�]r|[mV9D��g@�	�*S3�n�X7ڨP���Y�l�9
��b4O��9v�X��E�� ΄���J���u ��c����!Mie��4S���ȆJjV{�N���a҃����?a�c6���YS��Q���|����}�1�����SVv�����G��R/�G�ʈd�G����y��{���sĦ���ƛ�ܴ������\f^$g�="&G�Uq��������)If4`]��J���ٶ��ٖ�S?���e���i���?�F��X�jHP2�|���S���Ð���E�Z�tV���#���
�?'��XnZZ5��'�(��WV�0��]-0-���~�W洚Xt�����ٌ+b����Ee�a�7��D��1a�e��߄�
< ?��1%�.<��a��T��]��2V�~8�K(�����F������f:�-I����\��\v�W۽�C{-��H ��孽@�j�m���7:)��NGL�@�^�=���9\+O��M�\JO]M���.A�;|�h?�k2�ړ0�T.c"�F��N���]��/�1��&K�� �$u�V����Oϛc��箬:3Q���A��5�
��fl�!!��<��1ρX�c�\�Y�O�J��b_����y�_�)G;�-�:�r9&GZeU$��T>�>�5��O�S�����R�s��3��\N��Nߟ�w�9},�vёD��7˚��Ug�!��R�e=wd��z��0������]�r*5߭S��X/j�$q�����?�y�$]}ߝ�G�Ct�H�c�/���_Ë]�I��C��?>��8Ŧ9I��N9�}AP�Ԗ�����>ҽ/�A(HXj�i;gJ��ǧDKy�.�w��h���<p��v�q����m[�ѳق�.�-d��ᖹ�nb8x(��ƅQ|pT����&��Ǽ��-M�>B
�tS��2�v?QM3��x�ZZ�)�)�-�Ѫ�l-=�8./�4���y4��ʈd[Ֆ������>�'61��o"�]l��ҍ�5��_��;d�yN-=�+��.%�!�Ԑ0%���-(�#��UxTL}��\/�t&-�jI�m���j��Twp�^Z�����I�G��U}vĚ[z�Kwm];�8!D��UPb�>9����z�鷮�߇t��p��j+���z6��T�x-�D�Ó;'-wz� 's��+���}��a�FH7�!���	\�!�"0��휭�s$>�,Ҁ���j�����sc|�a�8^�����E�^y�� �mzQ�6���]B��>���!����Qch�Ѽ=���<�;IFZkS�q���h@�GN�x���w�|nl�H^�ȵ��t�O�� ����WYii��F��vx��-H�yO���-XT�;�=�����y�d�e�
�W ����Q�5'��d�^�ܗ6&�&	ꭄ\/R��W���ʈ�ٙ%��5���>uin-R�A:��S��2~v��&9o�����btP���G�������_D���h���),˘�F�$)��ߥ���_f���1�j�Īӝ^,y?)�l 3_9���dVtD7�I�+/�g�t���k�B�x�e���M�-�t=�|Y�W���Ը�A3(�S�*�Gwƪm"N�x#Li��o���M�@�K������������@����-Z�,uP&��ҞR��\��������`Y�oV�ۮ�&
�a���z�'���.�0�k�|��S�XѢ]���WH�ϋ<�2�|0���q�`}j�rH7���6�o���:鞰��Z{~�ڮnEB�� !��\y��QR_�N����phGM���D�|"�����1�1c�0��V�׻ �xG���~dʃl��H����6�+y��x�1���I���Ҥ���W�K*в��L�W�n��h�/�V8��+w �Q���H��_N>O}+�i#�\����A�;#� ��g��Ǜs6�M�N�5̘�ܼkQD��hr�(�oW�������j�e7�B}D�B$Z��I"p`$ו1�)*V����3]�A����ѳ��3�o^���}Y�A\5��V��{G��;γ �''t���S��W�A�B���q�������6�xQ|������y!��
��
i3����߈"���3�^$�J��S&���h��Ћ�.�� �C�N�7�,u���(-�/u#�R�x0�ՌnJiTu�x��,�~���"��!�:���d�;�B2����5��^����S#�0A�����pH�)�qn��6���N�ڈ>� �����]�B��l-���n��%�ŏ����~Q%,>*�&�To �W�"����4#�	�G��q���Xw0�����i���ھ���a�e�3S�y��?5�7����m$������9ۗa�����E�b'$$$�v`_%lc��|����1]�c�K�?�!�zd� ��&���S��\oF��
8�3� I	b*K�Cg���c+�C��(�_�o����C<��>�a{� �B����}Q�a���(�(%RR�,H��ҝ�ݱ�twI��ݩt���]K.,�y�������u��o�k�ĕ���ç�����&����Q�����c���:W�/]�3ٮ<Ȫ1B)�����4EAұ$��J��y�lE3��`���ŌK~U5:��۝�E��kWZ�h��`��Ν�z��]��Y3Zێ��j{_]�U��Wn�Z)&��ۺ8֯�ܖ��!�h�@�x ۭ��Z�_ݤE��Bo^��7�$�l__��N���g�����i��4�5��h��%��$ U�$_�Q���wO�+���c	�:�f-�-�l(��7u���D���u���p��{��ՎE���5�?�֥L�2�F!3Ah=��+��-�?�_��/�ܠ���<�'7�-%?R`���ܜ�b}y9�7� ��BFJ">l������Fi�Y�~zS�T�u���-��q]Z��t_��"a�Ӊ��d�24�fQ�<�-br����A%�.v[h��v�e��k���?W��ϘQ(�������`k�4�PV·�����hj��%4|��%��UB9�׷ߝ*A�-·J�ᬖ(ɪB�N�M�؈�w���7}L��Z���=gw*�M��W��/�|&d��M1��^ �0�2��bmAA������m�"�4E�Iʇ�r^��<M�Aj}3����g-�d"wbS���X���ù�t�J;���S�l�%ӫa��
��e� #G���#)'3��&���b��#�U�N�Q�����-:*%��(ƭ�6��s���� �-��ߦT��^f�f�,��-:�[�;"ʆ~`�Kxx�<~��k�7ߘq.ߩ�

*���~�MN�N���R:�>[��rNN�'�])Bĸ-G5�u~��/'Q$�@��7�Y.~��rrs�Q��5���u��� ��8��̛yF��e7���Ԝ8�b��-����pm��.�$Ĵ��D����9��]Xq��ƪ7/�|Օ�|AQ.iJ��n�Ķ8��"᱐f,ZF��G�֝����M�A�ʵw�;'����F)'�_/��uٝ��4��g����w1e)�K��3�h2UD}�˅��<�Ң�>�ǻ���U��
�f>�مtuoX��GK3�B^m����yȷsmo�.��:]Jyo�I�U�@��4�<�H]ΓY��۔�巙(rp�$<��qp�7?3��&��}ͨ��W�h���\��:�����?[YF�?���ۻ����A�ޘ�[E'�DA���]arK�f�������y��E��	��殭�7�~#�-%�����4�=�-	�	����W�4j�f��ik������26<�]��ׂ����`�4[1�w����TG�B����|�j�zu�[W��4�4"r�6s�-���jyy~� �#���[��*�nW����&WN� x%|4_� y�z����ή�ߜ���w����l�׃��z�o�n�].A����f���PU���䴢��"S����O��_і{��8�zv�7������w���=�ɅŤA^�"��A[ZyK77��2�����ό���.X���/�TG��{���j�#���	fŭ�T��W�AGl�����d�6Aګ��-���<���;s�?R��F��-)����c��Ovd�e*ˎJ^����k#ʌ1@�����ƭy��3mq��� MKZ��1�D���+�] 뛥�1Q#7+0�,���!lE�{#��y�,T��T�D@�+�V��s��V��
�kF?c��֮Ƣ4'c�~�����b�m�;����P�O��U�C��?��j�uY,2����Հ^vj��*���BȜ>娐� H���5��*��5[֣4N$$榾�K�AK\�?^�������>�$��+�!�첾��pp����<���
�-�|��<�`v!4�@��T!��(E�=�s����n��U��@<��ʞ�8����������?wk�S�ԟ�8��:ےZ��J�k�d|pUB��������$��*�8]`G�$�CԪU#m�<�i�嘘�o�P���Y���u�Gb��7���=�XM�/�߽vc�C9����d��{����^خ���$r�D��4�KIv�(�vkgCj�Ҩ뤚���D s'&�a&k�aQ����ΰ����@I�WTGbb"Q�D�Eڍ��!)�[�'-��0�LSU��E�W�)�qMm�TU�?jQ-�~:7�M���_xsD���4P}\u�����8}�L�5��O�b7��ҼBĞ	��*"T��컀�M����e~�5�ζ^��&��^����Ｖ�fýb]=^ !��?���0ѳ���_;�n���E�<x���+��f�uNN>C.�b'���C��
 �wE劊�Z��]�1�Y�WA�����3^%v�5g�V�s� ��W!ٝܢh�qK�9�u��n��.uzK�r��3ܤ�wC�i_��0[s�%�:��?_4�
<�){�	ҲBޕ/����b73C�e��-��Mx�?*I�7�)���<���,*`�Wڡ����iۓ��(�U�>��58��u�2�ږ�/ ��?�������9�W��చa|g5��c齯��\��I���~��Hfˌ��~V˖갸ϠS8_�KC�U�d���M��Z=�4Kq�"�u�,v�@Z�[��Dx�OfJm1��(	*7C�D�BH�M6:�YW���Q�G����^�4
thW��4�vA�_�j�P�,NU�=��d��5�F�o�F
��$���D���p�HQ�,��� ��;��NW﹪I�3�	**���ho�����RtC &\���Y�B''3`J��n3�`� p���Y�{���F����<�Cd�M��H�S������W8�%r2�*��6{^��%Q4�������Pr��;�B���lL��"�hu����GUބ|͹7j��0�Za؁E0�}q�RJ���M���T����ŷ�n����=���GQ	 �v�۬t�@�b����f�x�u��A�S֙�����,t~H������ 6�a�4���U�g��u�O�:!��wL�Jm��{��� yPY��5��v�
���S������_RH)��ir���)�k���h�"%���y��.�R��I��%�����_Y�c��u�1DP��Ƭl�v���H;���,�'�
6 �:_h�;�_N!��*�xX�1�|�N���.$���MV2�?\	�%εo8�=��G�7�M��	�f䎹j��>�)�N���BZ�t�:!c�Dͨ��gj�PqVu	bV��d����6)ߨ�X��&��X	�c5Ѹ*�J�B��5*U����i����x+  g��fJ}�{Pb�Ձ�J8S=�9�-�u�ʄ�9O+���B��������F��S�(%�hI�p����������$���\�~�΢J�����g4�o�P�)f^��
�srD��+�Ӌ3�e�|��ʊo�s�3������G�T�-�ApL��[ޣ+�3���dD4��BDNU㭧�;M��=���������,���"��doo�����H�����9���4W��J�ƅ�Q!A���=�Gͺ��Ly\3/g�̫9�+X�yJ��|��x����#�y�}�$2?ڡ%䝄�� ��%��"�H�P! x}�isV�۬|S*�*]��Q��ɫG�y����vb�&�1�X�
h��3~����ܵ��;2<JkS^�ٞ��tH����*]+}Ŕs��1;�fA<m�N6Z~!@hs�匶��9��#Q&<�����R�\۞rТ�:���,��V��H�!�����RC��#݄��Y���������Y������]���x�]�$[��l���_ ��5���)�Y�,���RQ�UBحU?��r!V~i*ٮ/ :����ޮ�0�E�w���ҭ��`߱1Z.q��~�w���f4��̌����N<�ϗ�y��j͞��P�d�-���΄�(�ǡ�kNFJ)1���˧��rV����%m��cPhL�#�7`jY��fA��0�1ּ|w�C�����39y}��e�9�5����g1j4 ՟�B�x�?��}��h��\Yy�"��˛mYw31��{����e�0���n����[K&e^)V��H�f�I�Pg�=�
��H�-|Ju"[* v���pn�@�~����7D��"����\� #D͊�}�q��? ��ԛ��V�Դ?����(n��ӿ47רI^T�a�X�	��{5g��}ۘ���-k���G9|J.�˖�j�J/)P� È� �Z����c�"*t��1���R�?�+[ɵ�����#�_ ��9�a>��>�'�s�n�*��zA٧���σg̌�$�,�q��5b������q���E���U�m|(��H=��ц�N�w�l�_Z�DU:D�vT�c�3+�[,�h�bB��Ӊ��������_��:��r���M��������L"����6}	���-�3H7A\X�� Q��i�Tj۔8Zs�yf���"	����v ��q�Uv�ԩCb��]DpK*:�\�R.�t��܌SS>՞띞Xi˚�ORz@�Ծ�{���[��ɻ�L0��L���Ov=vr�����m��{Z�3�x�^����$����?��H���w5d�K�V��[ۘ}����'d���ZȒ/��ʱ�Oq���a�_��ґ�`謬.u�������I��A�(�Ub���a�;-0)��Ȱ�5ɡA=�,Z!	���<4�j9Ұ{btc��H�n�u� QíAG�j��l;���<k~d	�}gMH�L���@c.}�멱<�����렋"��������H���:A�4�ڔ66��a$.���W�Ep�f؆M:��������/P1�T��J�BRv�X�N<�!{��#�oy�iyƛ��<��+�>��*���ނ��w]�=�ɼ?s���������B	�`�r��CJ� wy�:�1p��~3�N��~[��]㟋��S�)9�W�	��<?��D����b,Ʉ3RY?�=C.mCǼ�2����p���I�����0�m�e�)�V�J�Ars�h �֌����n����೟��<7���tguxd�ԭ�i�b�"����Pc�TuN�P2�����	i�\UHcl+sʝ��O��鬲����kv_��I�k���Y���4S3�_�?4JN�6��ë�-���V����'��BKv���~d|�;��
��`�w~�m��}Λx���/w�2��FI��:�(Kz�γ�����A\�=\[��ڨ�4 �)�?�����+h��\��Sp����੝٭ )�>t��s�����9���l��cs�LL4��1+7�����emYo	ص�ƓV�h'ly.�t~�3����QD�0]q�;6�֥l-�t'�f�A����1p�sM�}��ɒP8y�ǽϧ�rL��w�?I��J���x�V�s-��~�QB��m��F?7˔�mIK�+�������<��'�Vܞ3i��&�A�������N�ͱ�gć.P�5����Dbr��?
�f����!e�+t��G�D�wG��i�Ed�T��-4o�p?��xr����w����-���L�9���J@������͹J9���nK$��~��C̻�>`W nٙXD6��l��s�=��ħ��	l��q�G��oۂ��}��i�5��C���ZZ���c�k@~G���bX٘��!�q1���t��w
�*��uZ;�[�� G�^��Ϣ���F�]�r���0$�{>IL0i�|ZU�^J��{�	T�ȻLτI�%�{�94� � �tg:���?�+t-˶ܧMhhjO��L�~�l{��`c���Ґ��m$�$`3�06�񰠊���&H)MD�-�/�/=$�Q�8�W���CqHt[�jցW��6�8�T�9��z�{�:+�r�K<i?���}5��g�/ R'�
����]]#��z���dA&�G�õ/ �������Go���I�X�=r�~h� ��Y��s��qt���Ay�e]�Ί���4��s��j�Z�ԭF�'�9\J���֒��&��oi#��2�-��X�箥� uu��Dϲ�w"=3�5;V�?ŜJ!��絻������@�����[����|�A����9�,��ҽ`޿S��9���w�zĶ7�}E�3�:;z������X�l���?_��_v���Ȱ�� |n4��X,0�B�e��al�k[cx��R�)���cB�00iK�-il�w�=w���q|��E)E��`��Ү<[{��}]�:�b��#��8�O��:����s��Ϊ�x�������׽����A��PQ\���5�\��u.��VUG����a�	eiw��,��yK�#�TQ[٪�X�]-h$�_F�-��QV�y��8�uȝ�(I`)A�����!��E���fJD��`3���prֱ0Wb_<`�!����Ƈqi���R*6��G�^ �w�T0=��4��
��.�q�_��lԿ��'���LwaxO�����"��2����w�K!"D�HJ�ID'Ӂ1���/U��0-I,�*M��b���C��fK�h�3��d�9ɜ��$�*��;c4�La7��3��� ��ye��S{Ф�6�Н�~�$���:O�=�
Q�Ou^���G����%h�;$��Uc�1���Ok�Z��0-|�8��ު��+X�+�6��4��o���_经�Ґ��?����M�rȕ:<x�J���=ȥ)	�lΊ�Y  ���^�Z�bB����$�ަ�����߰Ǒ��K�!�%�PǓ�U�X�T��ÉOٶb�.L�� �e����	�W+��P��1(�b��TKJ�0U���V���0bA�HU0��9���w��D��"�d@ּ�i��ɭF����}Μ��#�P7�&/�PI�O�e�Q�ѲDeiV����N��B�ݍ���)�5��ܰJ����ɼ����:?pBjłT�$����3v�0-��K`�^�7tW�LF���kU�X$�Q)&��,>10+�t��T���o�����Lz��PJ�wr{���Jc��db�í#Ű ��������3'l+�R�Y)`�dYV��%�����<�x�d�ڦ"�[]������t���X�b8L�W��K(i<�y�F����YJ_'�,�45�MX�\�18����k�"w���~,;0ka I�+��%��  ����9��(L��mSk�/���I~'�XNz�̚"X+������BA����T�f}�6&Tm���zr�W�q�����Γ񺈖�L\�I��]���T����j�Ѻ�a�%�Q�s�-쫠�;o6\
��&&�3��!����r�R�Y�Q%��N��/�b��Kq�e�n5ΩFͪ�w���#�2>yE��E�%*��07��~��g� ���M�8�a�}x\A�8ض��zi#I"!�E�QMp����hC*�G�2�s8�gED�sA��p�"�
�~C|����d��c��zY"�����#���H<���߷��Lp�E-�6���X�h���Ĵ}�ԙ�?��b����wKL��`��A�d,s�o�iVo�bp���K��npo���n���}4�u,�keRY��Q�in��gb55�Xı��(kV>��q���m��a�`n��N2}�t�=����S��^�Z���61)�<l�.�s���k���X������L9�٠�S�D�nu�N?��IlV���H|9�����d�ף9҄�(//�/����6�%�����HikDC)��'����ޅ���ҿ]��Q��#ۂ�jw+/��O#L� ?��:�¥��Tq�/���<��d62Nv����WF o=�C��
��_%��� ��(�c���3q)�'%��<hԃ��#�w}6�Ae]~��:ɘ��a7/�ȝ餇��#�7�n-��7�0��2��Z'[KK���ߒ�udp���x�9��sz���u��e��L) :K��#r��v�����0���G�E�`ewe��r-�.\��PN�΋����6��l�.k\���a�`$^/�4$�ߛ3�� �V�ojS�'��O]�%)|�d*����ׄ�8.G�Z#}7�P�e�?!"���7�ϡ��	J�Oʑ��=��y�H��xy�%�����G�gp	��{+�qA��@�l��V>/�q��6�^ ���n�H����h�	��_������9�91�6v$�Zy�]YK�E[�����	��_�w��Q�gr�н�yn�3o*iD���o�����R������Z�g~$3���rj�/|��!�*�Py�]1�g��I�U8a�tϷ���<��g�∿d�N/���W��<�@;Cl7@����pڐߍ&>Rg�p����o���` [}�f�'����<�U���SV&���dÄ�?=�zu��^ �U�W��)��%t�O���;�5������?+-id��&S�K 
�\�����I�%�|E(�����B|$�}��Vk������Փ@r�~SA��U*1�LB�kR(�ҋ�z��bF�m�,�7l������a��׹��R���"w�_'MO�ߑ��R���I������[�6�}���f��f���8��6���c0O���5�(�T��ʆ%�%I^{�c��^]�4���۞em�	p�$@S��}��3m����{U�9,Ms�G��3_/��W��䴂ʵ3����q��p��g���2?���g�TO���^^(7	����@�~�8�����0M���@X�y�M�%%��w�0��RK���.eh+ۚ�Q砫K䢺~�����ߚ�sF�=��m�ᡨ4c~;i-���5�{�z.c�0'��"� ���  \?ےJ.���Ϯ��M�H�i��|M��`��R)%��3}2���O�7��b�e�ɷ��_ v$^aG�%�u0ϵٮ+>����exŜ��R-I�0ʝ�yO�i�Nj@��]�iC�:������Ą�X`ս�w!s�1D[ᣂ�2(/�5o�3�zO�eHR�k��]#?���\�#&��t����m�v/����`���S7���ds���m��29���v�5����bL>|8rZ�n��T���\ǜL l�:���Ą��?�7�Hݧ���D�3̘����mmͮ���uf<���#��v�n��{Ò5g�Z1� W�i�
c-Z��]
C��L��5g�3��r�lL��(�/�^UH���O�g�
XP=RC	�h�;@��2�^��HNР��C�e�H<�B ���sv7.����P&�5H^f�0���N]���z-D���o
ѢQ��j�z����T
#KEOs_ϥ*��U]#�w�I�6臶���qJ� ;3ʳ ���v�W���2�TJ����
%wO���M� ���S	(�6�o[9ywM��k>	
���jfJ[S�1y�3~���!��2�؛]w�����u �)��U��i
I����\/�4� x�$k�oE�?I�ԃ�L-�(&pC
%(�d��^�~2'�m�\Լ��JC�[���P^袠9��ٓ��{�4St�='����g}^iO:q��D/$n= ��*���ݗ�Ȗ��4����D�'��p�^D����U$�h�l���_�0�ZB�V�&��i��)��E�+��N��ʇK��>���Z��0kq���_ 9��'��é)g�V���>a�A ��.�'b�3]�T�������3�`neq5ޕ"�Z͑�v�_i�M╤�[�}��Rr��,���a�2 4f�����ҏE|Y8Ǹ69��A+��7n	�3p����d#樸]�������ePԑ;`����A�](�㿪�X�b^�JjM��u�kLR���������M��~%��_L'}� {���a������H��
Y#���������o]��Jr
�	�Ů��hޯ��,oq�d��F�s�f��d���{K�֘�ZZ�U�n�W�ejP�d�Ύ�l�o>!���[���Z���ؚ���fL�qja_(k�58��1)�t�n���� Ԏ��5U��LR;cn�IτG�
dB����Lȉm��ξ����J����uDbU�Z,���uIA�xK�`dSm[Z�V�_����\�]V\4��ec��Oi��,9�vMo{X��$��ǐf���Q�7&�z`��3�� Ys,��D�#�c�>�=}X�N&���m�d�3�L&aZ*�\"d962#�u(i<�b�𤣼�߳D(	��n=�ֳ��X��q�� ����|{�ڽv*��/���꾛؛���ڥ���H$0PT�J*��Å�VG�[���ۥ��ɪ�.��VC��Y�@p6Χ��d#���k?�ly��+)p$����uYD[����������i~�$�.��ʒ�Z��v��f|g��d|�{u��(�G�)�8����{��T�E��U��n*Ǜ�Uu8��{ʕ@h�o
��@���<�?�@�:/1��o�U,mMc ��ֿ7��20U.[� Ժ�k���핵�2��>(b[��"��\�I#��� ����)���@�%���D�T���C4	��6���Iǜ�ߙ߬@c����z�g���k@��Q�����LY��ǫ�q�\�սqUg3�ӬB�M@u�!�՗�c�=
��ݵ�ï+�Ś�3��\о+*� ���B9<�}�.�x@~�V�c"_k���Is��v�z�&]&�Lu7a(K�0�Rg��G��I�
�#BIn�[t�}��a. ��]�Co1�(
�O|�W��f֕�d�q]��y�b��% >F��?�(�z>U yc���F������u\�y�ڿ���?��BA��}kh�?+> ǡA�!�K�����}���1J�����vꧻ�˷�Ǎ-�N�%��$���AB��B6&��"��` ��?�La-M
��F ��J��𒿎5C	�'�I�1.P��#M�Nv����r{U�k7_8�ۂ:�0��T>q�m��F�kk�Hf[^��r��*�*��'���Sz=-m�2ޕ ��^xO�]˧ߟ���Z]��|
��<Ԃ��@a�v��/H|nD[ێ�T[[��A�����/���1c�$��^�9֝[L"^3�a3MCp/U��w�o{\�JyQC������ 6�'�����Y�,J�j1�1��(����@`V�ǡ�h�'wOD�i����r���E�?�?��]_ JP1a;���E�5�6W+ِ��>ꐴT&�E<V[�Eͥ� g��+Tʉb�>E	���>b��2 �v��Dy��	a'���Xv�Ӿ �m�ד;��3󘭇�VvRf��Gi4����v66�+`g:�Q��z.G�y��<�8�9�ͬ�~�L��)� �2Wa'N���o��WT�@j�8�W�q�A��?AH7R�_g�����zM]��Y�P��^T|�s����rEYHʹy��ۯ��֞}R������u��EP}�"$z������иn](J6��KpDd�`3�S�^�S=sTAFz.�PM2��W�gq��tnq��AŐ��q�(�`=?fn�z63��k��;��)Ga=Q�5}1ˏ��د^ �|jdZ���	^+�p0���Z������F�&�vxv��![�w[�do?T���N���W4q����5��GͱZ27m�U�*�#�*}�����U��c��`xݧ-վ���Eo3�QoҐ#��6�\h����}Xq�A��%5)��b�����3o��K�B��O��m��w�
L���Le|�y�����L�]խ���;�m|[��B��s�|���4˂C|�>+p��m���M�\u���M3��bJ�0W����Ӓ�������Zf$�^����*��w�j{(3'Ԍ�ӪNw��}�'.� ��>��T�k�3�n�����O� �}M������n{��c|zD�|��	$#A+��?m�V@�c�_ IFh��V~a~�n�"M|Y��hԠҿ�����h"�4�OG�=Ψ��fI�?	vYL�[3�E>�U������#�"��@�S�ٝh �H���L�夯hs�`��f�O-%͸��5+8�~�q"Dg`6GS��.Q�H�H)4��֢�|*���|O��5��~�������~nh�+�k�:�����$�9ʑ$0�'���e�����C�L�{�`�E���-��..+���p^^**��lE��tfi$h���Y��J�Д!��rܻ��2�������B� ED��i\H�4��;*���+��8�f�Eӗ����Ƽ_r����YJ3c��.��)Xlϭ��g2�&��2jf}L!s�D,��oY��26O?O��n�a`��_@�"�	]�f�wd߹(��<�PbF� � �����3@˂��v"PS�<obKn����[�Ȳ@����a 6x;�x��ul:�k��r�R硯�����f�Հ]I�8%P1��I`u V��(�̖��W�eUYQ�Z�1r���y��m^��ps_o�ʏ:�Ha}%�x��7���i�~���7/c�H��:�r܄���o~��dp��q��h{8ӓ�Ċ�3��Jj�rYƝY�����Ed+ր����D��ܬ���Qa�Fy?��TP�͉��r���������;o���	N�Z�p�^��J$�� �����d���[�j�@y�hr����נ���������|����>|w�W!��;���刿�.�����h�;�7�f���ρ�=�U$�4rtߥ@�P����2��{�����s�l�^W��>~�7�z�09���8G�ܕ@�ze��7����Yi�cƾ�D�����Q�9/�|�a^�~�Z�o+���u�b}��;�j7\qV�l���Q�A���C�GL�k�ΐ��C=��˲n����OYYAT% Ql�l_f��:9�d�UIнc^�59�{�~��sR���23����$����v๽)�Vccshm���D�]!�7��%Ъ�{��_��1�����a	e��þ]����(b��߶��M,��ԒP��
Hzb�������|&��9�%!�����R���"��1��i��[g޿�Y�]>�q���D��v��`�RAG
=�^׺
x�
�8[�W�+,�S��?�O�X���l���Z,A%�W����?&�f����;�W�n!B��Éُ��#(�B�W��C���y���H9��ƁG������+`D<N]�d1�L��)����o`{�9��{SUy�֔���[ i,�Z�`��2�Juf��b�O�ܝ�!������i�_��L�:I��#�ŲE�E��H�&xcT����U��$=��&���t���n��ڝ �v�l^���[���b �È>�bRr�l��|�D0��gWKA#��]�>L	�i�%�5&m ).��%�?��?s?�����=[�e�00r-�������6�j�Ƃ�{�U-h�T��^�)���G`pcY��{��s�k�ׅ�J��ʵ`yE��ӑ}u#x�`gұ��ɟ���
�{��4d�(Kj�=s}�5ppYv��B�t�[�<GY�28%��`aNFY�S�;E�l���3�w��S�FP��E���=����.�S��r7!;1�~�o����/k���
�J����S�N������J@MG>D�j��j˹�Ѧ���L��R��G�3P�7��6>_W�Sg;������W�B'd=L��2�1�+����W���c����/������y������p���i��qV1�fbd�-@5c��i@��A���[��z	'��ˏ\�êIQKu[>L�K���d���9v�Y6��|=�0�~q����u-�*uo�� Cj�I� �#�HI� /��ミ�q��J��~�Ķr����T���;X��C�7Z����Jj���C�.�쳮@/��j
�k� |�Csw�Ҿ����I��I���-��hZ^]z}!J�F�&�c4�v�2H�^	��:�/��4O�oN',ߌ��	䣌�υ\��v��Ո�S�.�D�o����0���p��p�0w�gcq���!H��8D���ue֣�r���v�H��ͥi�x~�l�����w;�4Z�1��ճ&����j}��np����9Y��	�ȡ�����n���S�{�$=�u�bDin��<i��e�1�H4w��w��b�FdO	N�bV��>��S�ݡ�����ő����[EK!C4��O^8�<T�.���2r�o�ٷ>�Y��6��>�,��=��-?�4WL�p�(�*� ��t�-�*�M(n����q���h������MZ��42Ý���4��S�*|K�1D'�S=՜����#5nj&���<'��Y﬎گY�WiIA˴@~$�T��61;X������+�1�!M��1���-�Ks�IK،y-�����t&���+��~U�u��K�pdg'��M��=�U5	���4_��ŜhV�HTDr�8UžPvN�G�"���� >����Ǹ��;M����f)�"����� �!�\AV���Ŀ�G����o(�����!��\� ���G��[�	��}T��ӊ;�{4wu����qf���E��`��`%aa�ǰѮ����7Ɗ�E�`�+���D�RTa1!��AA���V�`?�j���KU!_���)5[�Jei��2�uL+��F����gby��:y��C�ɏ���c��l�.�2�h�
�[����4���<� "�Wv�w�U{��L>���7�O�[FǏx~.9G���PǛ{C){}r�l�� ��*�Cu[�*�w�ҏ4$�����V��ͨZL#����]��b�����x��c�I"�Y�Z�ٚe�����3I���N�lK�������1ne��@�O�&Ŝe�T%��?���,�y8��]f��=�칫	������_�NG�ƛ�Q�`ᆞmeg[�Syc��<g��S��͏�T����1�+�c��~'[�K��V@�����^P���CaXy}}J��#˦n9�ܫ�����F��*_���E���`��G�OϤ��Q�Q@0#�j������v��q�x�'�_�\�u��
Hp䗅Ke3̍y��F�����qi�����7s<�ݝ�e��TI��9IBn�?�Θi��lS�uh�����ngb#��q{��rn�[��\�k+��8���V0����I��pF�Rw��S�>��J�.r��^�s־~���:7�St�����ח&�vm�ֿ�/�� LK�3��ߒŇ�V6�ܶ�h֞��N��|O]2�5�7ow�s�-������1�hN4A��mn~7.�D
�%��$犈
2|�[u������\�x����S�d׳]�4��rqa��=����(��(���z�����XČc�@R6�.���3��V��� ��^Q�*+F)e����[`�����m>�~�j�Ve^hJ�^���V����k������:�x��kM�*(8?S �x\<�Z�g0oKR�!��1�{'��K��X��l��3��X�Oj��5O��g�ivҲ����V�dEݻM�����ֻ�.���{6��mh�h�xͿQ��NRW��z��{Ǭ�+
E�m��<H��K�|����5F�{�)ex����q���(�b,�F��c�IT�������P��o�)h�\�m`9�T�p�,&zA������&b��J��E��@�U��t�t�E�R�`��_a��c�{��{k=�)3#��8��)h�M(:-��FTL�C�����9(�R�_c�2+����φ���bL��3%МI4׉�ϴڴ.m�e=�v������Ϊ�W�m�8�+s_M��TǱ�P�C %y�E���]mmeU���ۇ����us�#4�o@E��Ixg�	�<2������{Ǌq�B�_��ϩ�ó�:ZpR	0�{ȼV�x&3�ӳ�:�@��N�E=U���hh�fP�۸�����J��BJEQ��`��Ȭxx�G�af?I���%;o��r��K�YL��k����ٻX��%O�sBC%���nB�t��즫"�dN�w���#��B��t-z����q� eك�՚�.�b�9�k7���eO�8&,��!W��d����(JGU�릅��p�o
jj2�t���9���u{�fK��'�f��Vt�)�4w?�]��&�p+��fc��ǘR��Л����Vw�+������N��krQR��&�[�������ۛ�C��O���1!5�N�����M��	1V��zvL`�/B���9E�h�泄۽넺�iv$Re�k�0,l0�5+E��i��	]{T��T�����~��+����Se��0����X�tkn�E.s�y��ErV���ʮ(���ARPJZ`P������!��D�����C�!��B��������/q�=o�Zg�}ž����j���Tw�jG�]�υ7��)����	99Re��.��P3��[�T&fƐ�X̖0�rB�� w�ڬ�(r�Nd`q�\j}���\�3Xx(�����,2���+b��JU�I��e���E�s�Kc,<h���}M$��c����a"���ՠNQ�T@VO���q��٭ME�$+�|���9�C[N������O���������vi����Њ_���`�s�_Ęq<�}������@!�qU���d��[3{�������_L�!���N\aI�b"�#�1i�Z�.��?�H�![8K�/�v�<�S[ �������&�B�OH�è����ː��!D5{)II=#�Ң��T0��6��I�b���������|Z��[�/����M�ï�&�����tu��C��L�W��S�bf`�]���nn��rӂ���8�B� "�m>�Aa!^��G���E��\{ �P8�aJ�[����+�Q*W���_f� Z��h�կ�}!U���#QR/���=���='R��{#�����*�����s*^���2���r�hB�G����N&�*OW9ջ�A����
,I�)�K����n�������W�]�>�%9/�*��!|!#�w���;����o������$Y�Q�G��s�]e�a�����:�有�:�m=$*��K1=�ۇ�)J��Q8\�1�����=T�w���@����� ��6{vޛul�I�>��R����z��M��m��w%�J��h"V�G�'7���f��W����UB�^�hM�ߪYv"�9N^5N:}�4������)��җ���av�+��U��ڑ��D���������~�h~����K����y�6N_�*�Sd�4W�7;��$ ��k��BW�֮�|��VB(��_�����f�ŧ�1�\�h녦�PzMR����	z��<��ژ�af%��U�|8�'r�i5��+��
�5��`��F������հ\[��QP~A����?ǂ�I�R�J4�E*����m-��ֳ������?u2����5�{�;]9}���Lin�fK�`R�u�/���sο��l��3�\�7�}�-/-���5dn�Qtۉ�_c�f�x�K>��-ƼW׺BȸH�^t��5Ţa�k��wK����+WbNv����-G���m7V�݅����LNE}9
�^�0X	N5W�P���az�_�\Tц�QՏ��٢w�7sj�i ���05���,��[d
T���yĢx]��i�h8*�g9����
٤q���� ��>�}7I-%���t:�R ��r��U8����~6�26�]���6j���je�~O���];ǧ�NRF1`�-�^���l�z9�'��oS��bw�5mB�6���<�����c$�f�o�7�����e�~�8}�ε�20an��:z�I��vx�j�n��h�6.�7��[Fd�����~��,谝�<���2_R�fP�	 鿀�+�����y�>;�g�$�&��q���E�xNP6}]�`I��(��8�h�%b��v)�7��8q[�${��$>�|�G�.�b�V �o�%��Z�Kt�-z��_�W��rL�|\|9 �`�x��-��aSœ
�g���n���������4�M��m�����Н\�{nED�e�����O����
�C\(4��*��|a��Ӷ�kFpIm��M��4&vD  W �q��Z��>W����w�R���;��]Vw_�iIK��|j-/G��*���N�MĆ:X�E0����d��>g�H�ms9~D��	ac�
�ģg߹9ȍ7Mr����ӏ`@ɤ#�|9�0��D�kO�.�3�T��j
�i��A�:s���G��|i�5��#ח���q�� �dψ�x�_6�0(	���o�q��G��`��fAp���J�7١a�_�0�k�8O�_0��t���yn�֝����U�ֽ���mW�WD.=��^!'$��D����r*��7�ml��=�ӧ������>(�)��s�k���4H��,�
.��2'�	��_��t!;x��5�H��/�ju�R�l����UUt,�9�c�U�h�q��>۬�I �g��v���,��������6������֦��̑RW3,/�Q�͚$�V���ud��&صQ������! ��d;68��gR�O�:{F��ƪ��G��V.��Ue~�I,��[�I�9�֫YU2��B�bb�����-�j���=�H�[w.���=�P�oG #z���%����q�����ec�!����g9���g����' ����E�m���ܸ�7���^���?l$�>���H6fS���F�՝����e�<=�3�藽�R�T̐)�^�HM��)��v�Wk/"Q����a���.7)��6amgZ���l�5 $�߹��.�ʆ9�:Ķ�:�+w�̺���V�������6L�W�UA��N�jfE&t��y��2�5��M�.D�^yp��Q�Vm�Km�cPi|u|֯ϵB5�O�(h�V9��J�T��q�uxQ�w�f��q���%:�;��~{�dE��Zj��?S��\�qit1s����^��NS���BE�J�m��k�Up��:���bM�.��U$�ejn�Q�{���ℕ���j����6T�5�`�M�_\*��&Hκ��Ad����b%QcY��F������& ޺�5g
�k���$z���[��.�=�~�k�D�u�n��e�-�,H<yE�����)�m�́����'����e�����>���'���E�,�f����Kt_���	n��"Ct�)�`7'�oR�Y�F��ҨF��1̡Uc��#��qݫ�^�M���0��<t���f��3y��0'�M��|\�X�i�Ө���t8�-��O�z���Oz|�[Jw2!rA�E��`���/��?���	4��(9^�?���0��xܒz��9��|}�^���Eӷ�	���@Z���a��D���Z�`K�����}
>�7��꠩����>!|�tt̵QM�܊��o�c���_����~��:&���"C�R��(<?�u�)�s�'��K1�d�̴̪�r~�z��׍y����6���bY��~�Ʈ)-���plYx_9'�+�}B[��+%������č����a�+�z�l�2�7%���<����Z�U�Y��1	'	��;}9��O�fsc4��P�41f!��77���ٟ��[�#�!�N�sv��V��ќ-M��O��q��bc��O���A�\J�f��s�ܖ]���'�	��˲;o���	R/�N4�V���^�!eDn�sK@�E׾i�j��Ɂ�(_���j�4Y��ž����T�e44�|���˿<��G>7277XwC��3&����
�툭|��]��P��\�M���J�:��J��L������/K
kYI�.�Pl��\q��^t�m��_E�1�m���_¹�	��M^F�rh�ѽ���;^�Ū�1�8�o!c�p��2�-U���l��S��p��%Dfx����b�gf@��5��+��� Ϲ����KUEZ$�����Ϧy�,*)'���^c�Rkm}%�#��B��\�����w ��Y�r8�O����R�jǶ����Z[�*��j�#�}�? ���������a����	C��5a9�'����+3��n_܋$��R�h8K��M�iw��Oŷ��}�A�!�1n ]��$ �>�.�>�3�)�
w"N��9Rڜ�Q�{̕�Q�뽬��)'� ͸7�_�^���2#��{��وio�M����Ɂ\�W�O-N�d�����"2Z~���'TMH�w:�Q��. �����Gk�j>�IshҽW�yo�A�T��6��{_�	@r��.X���3��*^���5���<� 3�9eQ�����������,.�hK�
�	Vm�"���w�"���ɸ c:z�GhY��T���`�:�R�|�}\��A�8l���[ˋ� ���t~��It�-�ʸ͠�vi8����6��zho�
��n��VXT�|[R�����gR�e'y`tzg��bs��;M$�|"9rR-�����?O�b���]����-h˽��h
�{G�2�A���wz%�k�9��=�x��xi�O�$Ǩ��gz�̞��*$�� �^܀|��d�L�t6��ŢL�,5C�^<�1uB���tweu9�Naݔ�c�H�:;ʔƔ�>7��ۘf�R:N��T<@�PXI��F�J֫�0n��GmV�J�wt��B�yG��q}�\yw��+.{:��~����9lv��T���eY�ꅒRR<=���w=��{%,z�
s�(:(��ڣ1���D��5��D��`~m:"��7�y$uB,r�H�f��+�69�������i� x7lB��M��`�����v��ED��W�E�<�)��a��VV�����7���<N�`�����\ {�<��^~�QYf��֡�Ǯ�q��o�ʗ\%�{J��/���l��$[�0=�ؓ�����~�Y�k^E�ɍ���\��%�����-o?���G\�������`�&ho峓�&<Z$i��ՌQ�'Z܇K)vJ�s��-U�3�[x��bI�����m����{Ɠz"i, �Z��%�i*�`H�Z��ٹ�< m/YV�ul��nY"=����fw�v��8/�"��&�=_�-��E��|?�*�0=�`D����k���	t��(� [:ݕ�ќ�>$Jɇ?�Ғo�`�E[.�*���%��0��޶t�	;speǛ:j<U�:p�ыޢߊ�s~�L&�-	��`���w������ \f��`0+
jA��`��M������_�ϖ&[j&�密���=�t7�T0s����#�l}�|���[��)
<?��c�rb��-����6�X�����>Dv���A�6�O9�?�Z #�`e��������Cm� ���G<���' 9-���m�x����͈�������o��ݏ�� O����D�\X_�����q�@�cA��|���X���^���m�SE/�KܶA��>[ �e��g*Ni�*�BK�&�z6=.��f��J7o"w6�}����-�?��W{�,�7Aⶎvk�-PC08�-�x�b߷���IJ_$����TʼK��R��Kq�_��ޙ�R�1Ǯ�*��:#I�{ue���YO���]��q��xңKM5� V\8!��Q���~0�s����o�$� /=rK���V�ft�va�^�m+Q�,"�5�O"������ff҇'a���h��e�7��J���
��x��흌�T��ȗ����oi�0M��u� �*���@B�Xa��t� ��:+�����*�3�S�v�%2 ٴ��M%�˓L��뾾���x�Z�<z��*�5�d��A�����0��:|��sTa`"�lш�6h|���xq}b�������qu����8�$����ܹ|x����H�m5��Ďfrx���Fg��wܠ�y��e]n�����w�beV(�dObUAB���L�JZ��}9��U�hk��%̥t�k�i2��h�����Z64��f;=�����_g2�i���)τ��0ڻl~�:h1�v�u��Lp�!�9��w:��G�ҭk�lU�갣*D��>M��1�?$�Ǟ�S�xM<?�e ��Cg�/%�^�҄Q�x$C��4/X�`2)���1�0FJ��`�M��R`��fV�od��]�E"�,-�sh�꿫..Iw/�n)}Q�?�˅�7�V����yj+�	I�M��o��i�����!_0d���W�}�� ���I��[d��ڵU�ʾ���{<��[:P�O=1�.^9���F��3��Q���/���Z{�`�S�Љ��{���(��O���@�3��Q�ԓ�6�q-�|ĵ	M�U�>�ZI'(�'Ш���m����t�y�C�s�VZ�V�K��"P��oh�-gYߏ��z�{�Gnݾ��¨�������|wx��vq^)��L|*hL�v溽F��v�>�����^X��Λ�Ɍ:�3�aK�m㕴B5�w��b��k�_��:;3^=�����)K��
����y�MnX�(�2v�Z�W�T�j�:(Y7~�s�,k�뷌� ON�Ή��'x���U�NF���8B����ڲ}$3� �.9�#����`:j�o���2=�
��מ����GFI[3�i��B�L����zS��'�_A�E>�n�'NrֺR���u"n��̊V`b��wdHu١e']���5�N�|�`�Ͼ���3"rGі��p������8`��M�y���(KS�wG�ף���f1젂���^�GM� �� ��v��g/X�)���:��%k�A71�l�(:yN�����x�/��;r����ʓ�Y;?Z�9v!���ȃZ�>:�	 x ��&9J����!ur�͡���_3��?��ϪF&�#�a�8N��ޱ�Ϗ$9�D<�W�v�m���乳9�U��� <1�M#r���m�Ë\����f�|]�NO�����*��L�k0�Ga���c�`;kC:�^�.c��O!�8pǴr� ��0��㶦HS�
	�U/.�Y���Q��[aLT��k�L݈�imi�X17-F�uL��AqΏC֏��V�A]m����V�N:Eon޸�'x{D�j�����l�)o�ݠ�k����Q�j�d�#���[��/M��Rˌ�O���*�J�����R0�d���C����Fe�2�؀�pY�b���8�-�������2��C*�q��
�-�G�p�T�hEU�_����D���Q(o��nٷL|���]^�M�tt�ɥ���`��	�_�[�;ʴ;�/|�]E�#���:��w�.YƑt����_OR��c�|�by]ە���3iI���)���y�ZeW�v4�uZ0 ������g(�5��/?��"�r�����B��U&|���H�z[��?*�%{I�����^�}9�{���WU'6����*N{2��$^HxhZZ�w�.g�A�Nm�g?ۮ��!zu)IE�����P�QY+� �����.u�������.���o��d�ZYY���Qk��� �!&gZ�:�ވ�O���W��v!!�G�="�����K�T�u���d�ʚh?����Zc��o.G�%�uTΏ_�����|o�<`M\�.f��{:��;@dR��L���½81�^5 W�89g��;�³7�:E��~�-�ݒ{�q�1�m0��p��?I���n[��;��N)Ѱ��5#�/w�L2%x��'嵞��B/ߨ�I'1�hW^�}F9V�xy�|;�}����{�mE�ٯ����f7�B���B�@N�1��^Ы��fT��;Sd�-�lݯ6ɠ�.؎�)�c՘d���� #ᦗ΍^���ˠ����l��v�S8��G(��W�>����J��3�chڛ���Τ!E,�}}����D���)��މ�e�q�5�;Ҝ�	?
dȲ���)��2�\e;���$���/Fyܤ�㸺<�R����L/У/	� �
E$v��M��S}wJ�	�x����Uv��#�t�K񁮒��N�D���t$#�������8�H�������fM�ΰ�|�w�8��lmD�L+�ح��:I�f�!��=4�yN�	_��~�ǆ��Ƙ����N	�Oh��D6���gk���^�n!��H�W��)������w/jh �c�
�R�B�1�WWs3{r=V�i�b�$P�߉�(�L��Ϸ9����+�/��f���q����f�rk+�Z7p*���EX�VF�R۸�tg�$S�+g�[0S��>�AP�*����C��7�odW�D���=�	˯��E���RQ�O�H��O�kzY�
�{�����3��P������ϋ͟ �H����F"!���E�F�����^�!ϡi̇��rH��������"���������l]+i�W��KM���џ��\No�猼>�Y�EH�����C�>�K�̺o��w8�dz��wʹ������7���)�I0�(��3�09�x�x�ߚ�յ�RN!����ly)������	�緺
#AzF/ޚ/9Y�v���T��U�YDYH��XOV���#���H��G��uvv�����"^ƃ�!5V��FH@���������QP�l�Z�;G\�DN ��߂*���R����lo�Yq�0+a��N5�c҂x�ˏ'���.��t̢DL�iQ(Xi���~N�K!	v����=���MD�{N˜9ю������;ܘ��?ݸł��=`SU�h�¿E!��F�(�5׋;�.�ܗ�S�M͔�b9�w9������yAnSvIg�����P-D}�`�L"�H�7W�J�ttǼ�b=��>��ں�v�Wۈ�W�
�~�=˸#�E�i>n �w%���"J�a����8Y�nL���v嚽�kf����H��6���)�1i�l�^��Mh|���(����<�G�8ҩ��VH�*����N���d�f��9��{�>�䛵��U�� ���af�By�� ��:�r�u�����_��x�%8�W�-S���J�?�d��%l�\er�J�,�4��wB9��N0�+s1F��(ڻC�U��'g����S��Y����8u��r���ZM�B�� @m(T��V-赃>H��9�W�5���q�'6�G�h
ґ���*a[3�A*okj��h���ku�ȴ��)�A�Q���H�>0��h�Ӈ3>�Vɳ�mJ�	�����'��;ǂ����{��������nݗ/�<n~��yg���+�C�4��i憑�j��ݾ.�2�B�|x�e��P珩]P����i�O1v�Ͻ\�?��#,�d�!p�Đ`y3?^䷂-ӵq;�5c}�y���NO���ye|biz(;pr���vV��]���q�y�쪑gC<�:L��s��$
�f$VR?q���[?da'`�����0��\zEZZT�
�7�z�^K0s�,;�)����dQH�2�/�N53KJ+�n�����R�"9W"��S�� ҄�")/���4��&IQ�
�_ۘȽ�u�<w������E
z�$���8����d^x8d7���ఓ�#.h����o=fQ�˞�)���!@UD�S��V��~X�[ �������q`q��[����Ģ~rr<8��#`������֭c�NewhFS~]�QIQ���~�uc��9^[�G���Pe}�l%jRf�55��{Ƕ2�$��p�Y吨J�@�?M�R�Y!��������[D/RLr���69sT�
>X���҄SD��N�V�SL�]9A�nn�����v��������˨���d�3�,�͹T�E�������sg3Dxa�72��t4�D_&�A�t.�� ���p�"O4�g��#��\%C659˘fl��*o���Gj�r�z�����c��R�Yv��{���A��J1$�z�f����Ȍb{<��i[����ze;�<����
TV>1�dV�U�+�h&[�o�^���CK�I���׋�g��D̨���O��'�����]O ���{b����۳�E��'�q�P��	s�U��~�j$e �MGr��LG�T��id�]��v��?�I�4���͗z�KI��q\OT�	b�����о����QdC���}Z��#��B\���ag��s�Ǵ����Ri�ڪ�X=����t�EnM`�Hm�+�{6��L�hC!�T�.(����v�*�𡦐x&�x����>��!J3���)lq��ZjW0: �*������Y�)��������C<0 ����4���,;�r�ʵ�B��⡳��O p�x|��99ldO ���m�N�� `L��t���b��z���8ڠ�=ћQ|��1\�ķa�,|��H ��y �	-Mi�H������V�g�
H���p�dS9K�|�JM��3�Jk�P/�ݙ-"*�,�o��)�Ub#���Q��)(�>��':Չ0(+�.jPи�cB�m��V>�֬��sZ�U�v��>S$�]�`�]�{�w�<�����
J������j|��O��2�<������s\��A�F��]?�P�B�$e�F_kt'����Ͻ޺,F}��~Q_�'<x�8'���*$oj��f��Ŭ�o�e"���GS�Jh��J
�@�nޑ�O�Z�7c�ϴߝZU����2V�fg*�xUZ��t26�5�j/�lB����� Aa/�*r�R���֮_C����e��B�㸷k���hЃ�^s�MJm��d�}m��:vQ�;���DI�o�������Q�q��V��MWK)��b���Pe�{��X�.<��~ο���tU��L]�I��EI���o�S	�L��o|J�G���\*��	�Qn$?&S�&�����9���%�ʐ�*�O��q��g�wpք��ŖWVe��0�f��ݫL�ࣥ~�"u�c��Q���O���o���L��a����|��~�_4�*�Q�g���[-}p���kj�p,�	�) �o�N�WsXַL"`#8v�@�}��'F�+����+|p�FZr�Rx��p��o�������<M�_�o41%ϋ
D�����?kϨ��l���I����G���'�г8�p7��UFBZf��S�<�N��.��Ma�9�[��D6��fS
�e"푌�2[��si���l�HcW�'��6���p����pla����1$aY�y͋�RTeqe~�-�u���'g}��=�cv��㹺��#+~c��`ٵ�q�]�،���+d�w����/G�y��l�Q�jR@L��oQg��+�wu�)�Lq���3m��G(H�=�Ƶ��f�\����t�Z(n
����i�(q�uvR�1�rUޔ؆����9 z�@�B]�WM����N���K5~c TY�G�f����\�хzټe�-�)D�`���g����Q[3xh@�a���ok-�E}V��l��"X�b�k����[x�	Fl�R�;,����t��;��I�#i�=��Iy�h�_��GRR���Q`Y�t֍WsI۲=�<H��sMx�h�Qf݉ns���#B�G�M�{4@�ȓ�z𦻨ׁ9 �k!T��I@������<�y��(�9T>^��rS8�F�]l���9���Ww�X;s�e�gӻm8�����V��ϐD (��,���eqMa��p5����SD���?EI9X�hp_��E�	��/�U��n'u���H����b�XOU-����s��H)ZE�
��0ku�z4�V���0a
�H `Ԫ`j
���s}}��/�P�ݏFm�P(F��c_{�r�q��=h�>י�%�.f	����~�'�C_IƢB�v�G<�xlB��UU@:�����d�ծ�����d�l�cÒ�dY�ݮϧ��=$��4�?K�G����S�i����u����`,V���S����bv��r�(A(���|��G��pB�"�� "`���r�4P��{:���3_�OS��#��ʿ��� Rx��Е���%���}�[��ʠ�g��e���]ݮ�!S8�f�_H�W�����5V�<d�5?�xqj"�֦P�t����ږ�R7�;B"|df�oG�1G��F�{}�V�����Q&]Fb�v2!�(��������X$���I�g�#8���w��u2nfǈV�t�5�ކ�79 '�.���t�/�tj�|X���w*�܃i�H�R��+��ʗVirJd��Qk>x3ּ_��}��j�9>��>��|����!/ϣ9+��S8q����v��g�z�'�{�mK,��\���^����R����i�r�a�A�b�<h�x�MmtRH�im�$���D�a��<�wD��\Ɯ��f�#��p��6��BL�sw��ֳ:&��3���l���	�nb�O��_� �Q�ah(#/G��`�8tH�cJ��q,�E�}C��1���+���(R������'��٪��N�3��	�A�_T/�����HkKu
��/찮@�Ϳc�v@R�Wr6�mnU���z�u�Q����f�[`*�vU�����]�ǔ�G��cI�p.���PNX(�g��%!k����@ܹ��R��+5Cq�2����4���5ߞ`Bw� ���++��v�S�*c����a��9���qY}eB`���� \.�Qī߱�V�N]�;U����>KU>jz�_^���s��_Y΄w��ȭ���j�)U8ɢgy*P�n���)�:oc�,�5m�7B�Tgm��ZJhN0\���фu�A���q8`�i4�z���.w�ǖ���{�}�Y�_U�'��t<+
ǉǖɥAn�K�?�<���,�8аf�^<(�'�9uh+pX�*��N�7|�J>���I�򚲲����kM��n�)���q��/��1�enc%����ں���^Gs��c���x{��̻�Z[q�ɕ�msAa�Qgp�����Z��$h��z�c/Qn���f%X!\��a��>Ej��|A��<�B*���#i)��vJ�41�¶�Hgݾ/��rqt���(�.Ԍ�Rp��!̊�$�LcȨ�b�.n�=�*l�.��J�:�s�C�狓u���b�|$N�^�H�l/��dlY((�sP�h�h���a�s ����ס�����m�T��1U�B����Ҥ͐�2K��x�5LK9�k���,��#C@���'�\B��G=b��VM�{%��>8�}�(�9��Y4C��պ�>��7}Xz�~I�1������砂�#����z3]%�u� ���=x�z�����H����sE'R�寤B�$��`��_�I�P�k.�*�4z;���}>n�����E�mq��[dU�	ń�:� )�5��<Z>�������HM0�5wd�!��?���uew,U�w��n�^ĩg	]�]W���?��55M@��K�w&��rm;\v?y�~}�Y��_���}�rD	�ݴ�ݏt[Kqƴ(��̃�T���L0��!/��op֎ܚ�]���0�KPIJM�^�F�d[�N�rXO?����x�\P8>U*�a`�Xh!��ݝ�Q��ScU���`��O.	�P<[���K�Ɠlꃋ��>*�a:�!>O �©�7�#��W>��Mo;6����Aŏ�����PuͿ8����q�u�Dk)/�ݫɾ,=v����8�T�8�k;Oyky^tP���)��m�r[f V��_R���ha�ݽ��4�wɴ�� ����{�ƪ�@, ��Ɵ�����n�ca!Xk͑���t�׸~�����]E�ɕ=ɋ���K�`�����A�过����d��G�b.pt�@۹����=�E5���DZ�-.�/Y�aSפ�@5���J39\=�ٮgΌ�[_1�m�}�3��� D���f���<,4�1d������o0�g���QT%XD��R��P��s���{Y��TA>K�����\�5h~��2��"Q�>ZiqD�.]�u�xs�;fO���S쵋���$(��`6/��Mr_k��~<����5nh��-��K�����2�_�֪ɕ�T*��KN=L�cho�1i�P� h�&�e�Q��������hZ5��8�d��׹��*_@w�і�s������l/B�Wt�e�j��!���������/�E�m���p�0�T�v��二r/��+1���p3{��ځB��4&��j^���n�o���#Q�i�_^��'H�T���η��??����0�$�#}��ӻ����ݹ�f�B\MF������Ԅξ�n�Fv�#��� �ᓻ�����yo�2i��JcYKͳ��B�����_�xO ��׆_r�=V�dˬB=%���ŭ.޾W���>�3�>�$��-�o��EE�o�]�V�T&�Pq+�1�Z�+�I��@��|r��]¬��Ѿ�B��(�;��k�kX��a
9U��$��#Ĳ� 3��{���6��$ݘ����?�x;
	V+;����i]�&(S�/P�x�m˼��`䲅���!�t"����@!^t�Y�	c'EDC[���xJ���_�E4 �0g�q4d�� <rK�.��nE`�ח��ې>�q��^�S�
��F`�����)r(�Eڱ@p�"�P;9G��K7����<�>"��^�����*x�w�r�:y:�9{��L#x�Q�>'�-͆J_q�����Mԕe7�����J�@KJ�5����>'!�]f��pđa��)�1��G�ޞ�.	�2�v5ozf�����߾7}f��R���ڨEG��;+K>JU��u��
�{�@��'�5��z���Ŏ��z��+cF��\*�.�R�k�U~ �����^6�?�y�����;����J�;�"ݶ���"r�%��w��8|�%eB�aq�|�uz̋6��]��?	�a��B��Vk��7W��u.�wY��f�����_�ƕ��쥃�n��t�F��b���t+��i�r�:�g�����"u1���%������*|d���lx��wOϺ�����rE��}�<"Yv���w�v�$��Z��G���t#��b5�y��P���mU"��1!�;��,k�k��v�r��q3\3�{����_�Xm6r�2,�e�굫׃�t
������q��U�j�=l�:U.�g^�gn�8͉M/�G
��ނ�+�CE���X]�勚o�;��z�^���2Z�S
�3=�2Q�l���l��ݾKx��K@�n�HT���ꉮ*��p�u���
?Kz����P��D]�W��Ʀ�s�S�HhǏZ��R�{�η9iE��#���t�b��v��ġ��:ςbi�������BO�"�R;��?�5T���f�AEC����d<��S���:�'��jO�:Ъ�:&M�	���<>�R;Y�Yyh��rA4��(>�Uj�g��9�^�9����)d'�4�v ����6�s�R6��T��x�B�_=�k���3��eY�]�ي����BAhO߇B�d �N���2���!7��<�<S���}[�l<wAE���G^�K��pܴ�tVWe={.�>ċ���H|F2r0A�Au&�@�=޽�}I(�U��H{�����	'(�e���w<�c��[�o�[����DJF$"?#��	���!�&,;�~�,ݟSU�ݽ��}{&��>�z���#1����`�tU����3�n�����v�?�
�@<�ŵ?UVV�עB/D��=���8lgq�=&wO�U�r�,8V>kOW��=w?�yt�:7{x�YZ����u�b�v����r�o�olG�R�J��?�I��O�1B��^N�ߙĴ��	0U�S:���OV+9_s��IGL/�۝
�R�4�8���z\�A�t�.���u�Fϼ'��߯N���^�?���_� �BL����������
&`�}[����uJry�kz��9+R�[K�޿�����`r�_�k,3�\8<�헇9�iQ��U6��)�M]<����N4⁜_�lX+7�t�m���n�c���C)E\^���*�fd�5�W�0���6aS���ގ�v���lbbuN��:���MZ�Ru!z[P�	����Z����"w��_�j$�o=l*R#�rJ��4�w����q����������ˡ�/�N�c /���
[��~G���{i���a7 �
���zuhJ�U�?�U(�ڳͪ,�9�X٩5���N�������ŸO���󩭼���~o�S��D֊�Z��GG&��5\�lД:%,��CVՅ�fK_�|c��^n��j:��*�V����Fƕ8�� �A�,����(7:Z}���U��_k䫑��IitcU�j?�5�Ʃ--Wѓ�`�ytH�Y���kd��O_��P�_�f�B�}�j�^D��|�{<��^�^W�g*�k��BSm�s���DS��A(�q��cB���M��{Xtq9ަx�R���O�X^���ݚ�0{
?|ܜ��jT�O1�]\��>����S"V5�Uk+����p)���cY��tGibȆ_R���;f�0s1Z��3���a��,k���G�Ί@Ы)7N\��h���`�wlJ��\c���8�!w�r7�Xҧ�lY�~���n��m�?6����{"<�����p6D���5c��U'�t�!N��s��L3�k%GXF��8JM�M#LZ_*�?����������KJi$F��R�%(��ҥ�0��N�DZ1	ɍ������'>��?]׹�}^��z�׹�}���J��v.�{��v�b��0���Ŗ��\3vWwuޯ9���J���PU��r�Q0i(����	�@�
�_!�N�Y�P�EK�����,�z� j�??2��#0SA�ɩ�vB�Y��3׶3?*F�Q�l:m�5%�9�e3�R��f�O-_e���~�W����q�/�4GF-��'<�s������voT��l-�3 �'�~��N��,��71f��{<9��-ŗ)��G"��>x�.��~���q�nC����n �ye^>m�lvF��� N?9��A2�64���~�o�1���˚�w���c2>3�6�>��x��Y��Z�(ĕ�(��>�������UſO�@�Ζm���_�ү�n��S-�1�q�-����m���o ��G�;3�>H�'��h	����(��K+P�����<�J�X��;%q�����'��Z�?\ġ4I!��/S�2�������)��=l�Z�[eQA��)S�ab˃�s���"=�����J2��TR��nt�.���6���-m���<�8���[����Yֶ�v�6��R�NC�!0؛���sbխdpN��ۧ�w�C���S��?��%	q��j�s� t�(����;']0ݨ��uS߀7h��0=��7sx����!�Yw��Z��5:����^�9�&'_���.+���_�	���"�;T}�L�*n ��x��"4<E�q]��r��U�x�H	E�i���v�����|R����%m>%�g��� �I%�
3E�gۃ�"J_Bk��R
�*�X��l���N���me��E�icb�Ω�L��������^Ε�L@	���+��U�rM=�|��X�n����E��K�F��#?�I�+#����c"5� �u��*�� K[�]Q\���}x��;([��T�/,�'H��v�1y��5����@ߥ�SɄ��e�+i|K��9ȬR�;^��wD*T(�>���f�|9�N���D����C?���7�s�a�� �IV���d��Y��2�ӫ�|��+;L��3}��à�7��Y"�c��_8�P���Ny9b�uC-gR����b��+<#�T|4��š�o�
ݾFK6�I��	�'DB��E��p���C�+�h��ؘ��E^U[��;�|p�Y�Z��疝C\d^���1�s��X�`���4���~ q~���!)������%W�q6��R1ET�
�OmVf�C&B-��e��]�$��װ��la�7� b�������#U,r�^�/�`�ܴ�&n'~r�U���yZ=M^�X35��v�w�~$��Ǜ�����/��k��b�uyAn���ڿ�}p%����*|��$s�� �âPԲ�t��u�}U,C�,�6��������4z�"��|����ۏ�� +��f	��o9���$
�[���@p�]`�[��'Sv���� Q��?��4��)RU�@z��J����v?Ɨ�>)���Sv��RD9;�{ꛒ����!4� ���~��	4�b����qN�b�VK��K��xqe��,�i�5,���(^�:��5��:�8A7x�r�O.<\�����5�\oAw��:��wW\�_l>�H��CP}q�Rb��ǃw��`�P�@�pN��C�Q�ǔ��o��;��]��o5��}	�Z�{��$��T^�R�t�����H�u�q|��5��@WE����Tl����ϣ�ݨ)P,0xyۡK�u���ѵ�ݖ�gb���-�̠Q�1�F9�βg�hFׄ���ܫ��V�?��>$P��Mk�c>����ˀ�H�{����wڰQAݝ�Ku.*�8��ۤ�M�U�Gl)�cp3�9� d�0�|�KE*�z*^��U4+����ULB����'~TM�%�@��CWE"�/���7�5?͐��6����i�����L+9"�8.�W�q�I3� Ќ��ن�fWvȫ�bU�=�%0�b�V����mE;������[�S3�uN�]�,I܃��U�B������}aH\�p��ܵ8�*"�ؓý�c��l��p���V�d7o �j�ǈ#���b���i��qgp��=���Av?c0�T(�Ţ�x��A�1,XPٌ'M�S#����
w����B�ٶ�m�ٕ�di�~��x��r 4Ӑ�$P��O};�g�kղ�M�pm�dEK�܋�Ʌ"���� )Ͳ� D�*ٞE����nw��4�����4Ġ���R��yJԯL7Yc����<�[8��;k��L\�c^���Qr�71B)c�
�}a97 ��֛�Τ�����,ͧ)���H�=ִiNkv�+fB�����k>���������i$�G�ci�Ɋ%�J���Ij������,;����)�0�p-Y��	�G ۼ�4��;����h�&�p5�NiI� �d���Y�Wk�4�x������Iz>?ƻF	��χ�����X�@��v~Ć`޽�G�0��>��^����o�H~?�E�w�5m�"�a\���Y�z 3Lmy���>�����!��:X�3)6��d�P1!��/y�� ���ш��;RȾ(����J	b	{�]�\k✋}¾b��8xw��~K	�Ĕ$є�"��Ԭ�e6� ���i-?�v�%��&-JY!4��4v��P՛��T3o5�������3}r$~��������O=��j�FX�=�f�,�1u�p�خ�J���zg��ؚ����~bq�yk>��'.��RZ�ٽ��p��oW���ͱc���2�B8Z�E�g�ot;��t[bRT)�>
/L^=��;-.U5	ɳ�D�;����ѥ��ɂ8�ڿX�<~<_��{),�oڲR�m�dO6���*���U����xS���@t��������粤w�������E�k��<}���B3��/4����i5�12q&�Q�S&�0ذ�.:�?(M-Mު�D����m$� /��A��� �+#�
w~ +b�r�J�q�"CÄ�)�4�v��ƒ����$���Mn�
K:<��x�N����Xb�!f���a�*���mCT�U����ߟ/�~l�J_�	 �A��NwS>����,���2xc���9�h˖�V���&(�T�w�+,�f���/����Q��vNVW���N�<�����{�C�+�������\fx�҅��רԠ�� ��I�9�v����Co�1#5��ԍ�E�~gl4! ��-Ti$���o�J���G�t�B�**�}@,�gt��4�J?���T\�٪q���!#�sg����M�f/ǯ�7�,�hc!��RN�X �-=��k��),V0�]�X�.T�J߲��*�hzg2�|�V.ྷ|E����� ϓd^c&'�7�9.N� ���i�N:��@�4�������K�߮��+D�����2�Kea�A5꓂�\��[�[�z�qph����>��)"���EWl����&f0����WR�&��l�Y�������7R�u�;����Zl]#�j�+k��Zʩ��F�$��sf0�`�vl� ;��FY/�"Ci�#k�}żҠ��;h,Q�$��I-��ꩤ��QI$��I���'�;/�H[�AN��<a�iAZ�+$**�
����ܦokW��ҺZ{�G�M�� ���aL�i/�����_Fހ"J��ޙ��%���ݱ��zk�#l5 Dzs�'�Jh���ŵC!�Er�T)����4Aj�$Br>\g{��M�����K ��)[KhN���>�d! N�J�<R_�PT�LÅ��7ǩ��${@�$HLwСT�wW���I�+(O}4��(g���f*��
��q�!ʣbO�k0|f���R&x2�Vx�����Q�8��_!Řo��R�:�OA�ih�%��e^��CB7:���C%�d�Z^��L�9�(�,0�:^Zͥ�d8�q!�jF�CT�����W1½A���X�r.o��r4�P�r���M�J�����!e����x�����[�Z���W��)�ؠ`���ˏh��vWz:�g�5��}�FT�"�W%'j`�㻞nyQГz;�̅��2|�;�ky���f� >�>M)ɸ3��!��xŵײ���+�2p��շ;s���j�0�۳�Z������������8���g�E�J$oQ1&9$3m����|P`�=R�/>c��v���Gϰ�5��蛾?��9��c��q�� m`1�	|��߱�X&���3�=Rةf���-��7e��	��\�؍o�)UF�ksPLA��ފ��{&'z7rb����{��N���T�?u�Nb�J�K�$�@5��4
��s�I��<�Ws$�a�ܠ/-~m��7����Ԣ�ˡ����0�Wo���o��`mJ�y�Lf���"D�s�}kJV#N��~�N0G��>�:�A�5+��z�V�nLd�rz��$
���@�iè햢�C�z�x����MF�>q���r���j�uS����@BOx��>�������w}oi��cxޏ�i�4Eh�qo��W��J����O��s���t�+��f����_�`�R<`LV�\�����B�e4�v��[ �ꦤ��qn�L֐�]��2�W]���\^�k/��pqzׯ��.�?}U~ � �LP m��6ۈ���[���>�|;�C2ԯ�7f���:� ��|�W��>,�t���Ϙ����*�h��̈́����?)��I<?X�<*=����*�?]y����K̷�.�{��jz�N}�K�7����W�6i��6�]�R���(-[#eo����n|v�	�AV���3yYXYgtG��<���o<&��En >Z�b��߽O��΂�8M^�Ljo�t:��
������:��P����ųj�U�`��K�K *>8՘4ڜM�u�Kч��`��H7�By޲�V���c�>Ɇ��>�x���c�/���m�,��աw��D����j�� ��Ϭc��ʱSڦ� b��'2!�ٍT�E���H[��n���;lƈ#�ֶ[Q��r_Q�J5��3�@�8R57�c�'۹!gL���D^Sr��a1iU��� T崎 `����I�%�n�!����O'P��%��;���5=�_��H�`�s��`(��1QnFS�:���F�Y"AQ���n.q����'�O9�(���K�%Kdy�I%%]�ߤ�`C�w�w)5�v�\ u�c�Z�@�X���s��YJ�}�0BUYK�{S�����n��D���B��$�9��2"(�¨�����|��#t������h�M ��,��t5�J��8�B��G����_#}�[�H?PzP�o`�Z���:�#s���`�ݳ�������Kd[�'�59Ds�i��iK�`�26�F,��,	�p%F�bϗN��5C�-=�8����p�L^��mn�Q>2x��F�/����"���o���5����ǆ�:D�l(���T$�ꊇ�W����^B*�:����K�ur�q8�Z���#GN�/�3ŎU�b7*��OBH�7؎r��X�N+û ������ڷ�11�p��|��E^FJ^~�2�U�C��p~:�r�Q�}
ɣ+a�&����e)�Ġ���O!E��c:Z��*K�A!Tx��4�\f�p�Z��od���3�Ls\!�L�*b����0nYK�!ؐ�UQ=Bo�_�9��l�[��/�Y�y�q���6��A0��l��)>�yd�	�d~��]BM��@J�U9>�[~JE��ܨ�K"ᣅA��{�ϸ^JE��_��{�nYds�;�������BAt\�Fe�u���4}�p��j��ڥ	hr�ʚYYK�I���m�����-�eQj����؜J4���.T�T�q��-P(�F���,-.	�d>_��Z{�K�����F
Eژ��7D%����-dC�L�];T?]��*�@���B�x���1Ә�Z��K�����:i�Ҍ�@0_U���z
�����h_�_�d��u�A���-��&�JDqqEc%@�k�YG���"M#ʽ5y��S#��H��*o��1��uQP\�*��d���py�16��a�)���^�O`�uv���2P��a�2~eۭ�֘'�hZ R]��#�7moir��. �.�H�f)�;���}��[�h�VN�=/rRb��M�~�>�g^�ldj��_�$�3=VvP�Gx�k.g��t����(�	G�/Hy|	��w�4�h���
���X�����u�I@��o��poy�R�g���z�w/uK��;�}iR�>}���S����Q�ߑڳ�ٻ�S)�ݥ��N{Pړ[G� �zݎ��o�MN}������������X�lii�Sk���;+�?�Q�F��c�sR��wU����Me���
o�ߢL{tb0�E�$�Z����5�ʞ ������ye�Eޛ/���n\y�*߷D���	�Ӽ"��H���J��5մ%D�3Sǡ;�jەKպ��6��|�t�W#�snR�K�(q�7��pR��-�����e�����5NcB�<G�+��AY��H��Ke�<�ƴ�����jEt<����E ;�n��;��ͥ��TG$J/�l��X�J2Tsx a��F-9W����E$W'}�Q���#�i[PGz�c���:�f����:�Ѷ�*����O�iߠ�zVEA��ύ9���|f��"�zbDэ�P��a7{��A�W���wt�\A�W��W���i'�"���\-8&s�d�,%_q�������0�WYKV@���ޮS��k/�h�J@��e!��α[� �� �ɧv�uwdϨ�YbFP� A���u#�*UV�ϝ/m�I*Y�����ZYt2�|�5G�UlS��Ua���N=ǌ@���nf��W>�,�͉nA,����r�WZ/�(�ܑ����n ��ca�L�hT�.��BO�~RN��8F,@����2DE����''"��2��D�&�1b^RQ����{�,�_�"~��~���B
�2\G������P=^9F�`ddN�(��LiLe���o�(W���� Nβ����=p~؀;�KO��l;�8Ё�loo�2�P�:qz�[��#o���-�C�C9&RG����U;
Z=>� a��D`a�����л���y��&A�9^��C6���� �V7����6��5G�g��j���Dfq�t�Y�
��\g�·���*���P��.�4H_�2b�PO��*�j�b�1S�񤿷w�����/���t.n |�� �A+!�(�����L"B;%;d��o�7x��Y� ��Ho85jq���`�kF�H�.+�{z�[����#�����1o��N��n��r����^�g���J��w.��1ꮜ$&��}��)���Yjy�}|?k��IH��2�4�z��a\��,(C���"h����U'4]��k�ĠT��m�Ll�3�R�����G����S���@��?~�������<:缸�vohGw
_}�`0d����<�����h*��]��Y��ݶ��b3fo=^���겑Pg"�j�%���������ݲ'�T�;��6�^0s���+^�g���3v2��Uۨ�_��?�g04�$�k�D����6�]�/u�NW���L�֮� oꏔ�#���G���VQ��T��=�Ku�K�u�ҧ�po�c$m�O�j�k3�׽�# �O�$t���L ����uZ�Oq@�"Ua-�W	6|.V�̜��8:��'TV.�h��zD��p�����'h�,[zݚ����
s��h�n�}�l�Y1��B��d�F��Qg�!&�������`�i&����5��@3�@��cic*5�5���⧒�f�0��pY��d����f1X�&�'C{{eʦ% EJG���Y�}�q
�q"6萌H4w��k�lBW�S!�> 1ir�+ʵ�s\��1�l{_���_x
�}��r�=������C�MJ��Ay�5�$����*��-�^��LJ���-����Ӝޓ֞RllDe�,�TSn�?	z�������3\��ǵ���ʛ��$�AESk�����v��y?�`�v+,�� 9�b���f��4��|���o� ���3q|z�L�e������[ҕ�~>�����T�6��ͧ�)��O�޳�?�6/[Rtk�z��VZf�4L/m�jX���@�Jŭ$�S�%L��>�a�DP��7c��q�����,��ػ�~���ԧa��ɛ(Y"�mk3$#�]��ً���תjo�~�~���J��P�m����/]�~}t�-9N��w�`a+ї��}5i��M��?��~2���d6|t�
�	�E=>5�5�����8L��y<��4=�c}�i�5�y
8���Sڞ�!i�G	dNfW��������P�)n]n�(�K��\��iC�iʄ��	���2Y���Q0-M� /t,[!H~� �xPOi��m��e�<��a���� w~����g	�����<O(Q@||���ط��T��d������a�sQ�/`��2REpg2�k���J��OzQ�a���Đ���f�+�1�&���+�^�iHWM�_��a�_������F�����JD�y��~%�| IzA���ceܬ"�[p�`4[�B�����9W�B��H`��^�?M�G�������N �Fյf���;r)=z�\��%�s�~���«a�Ե1�b<�$�9��fuQ��_����˝��fq	�^����@7Ug���|����*�S�ep3|U���?r��������P��y�~�ذ?�a�.��g��6;�f<I[5���-��";}lT���z�Be����fPc瓰��i�A�$)M�f�p?֯4αx�T0��~��駶1:ǨrQ럻�A}�;x��=���m�Wk�(����Y�՚Վ���,��S�	���7�S"��g[����K�f�x�Nk��t����m�Qo��à	��΍N�Å#�ٙ`�	C�+��&L�E3^���.��废�L_|N�_�4WL$�ӣG!�[V]-fAÊe<Ë�?K���\�c+F���W�Z�]�J��>ـ��i�HQ٘ߞ��I�p�z�uR�éNAɬ2FQ*��*��d����%����Zվ(W�
�!���:Y�^eV��낁�;��U[���{j*�g]����_\W���.�i�����j-=�	��C�+d�rܽS���N�E+f�z٨u/6�ii}��ª���%�ݵ&�J6}MZy����3����?ؾN�"�)V>��0D<�O���q�*r�~�e�y8�NM�I���^4F��2g:����-����|Lx�nӴoג��k+E�>T����mk�P��]�gy���}����3YX�DaY!~/��H����˅��ݯK���>e�yJ�A����o6�������;�Ϲ]�k����-��K�΁��ɇ;��.	P�̳�Ƶ���ow���~�\d^��/��<��:�@�,Lx�]؊N=Z~5��ЕF��"S�D~�.��/
̸��M�����<�i�?\����j�_��G+���������2AP�3G��\�)�à��v����]���J%[j%�\��T�S���;�������x�b���^����?A�ƻ�����&��
�i(ǇH�R��2��͜:J��j���GO3+H٩�>�_>��9�}�K�U�������]<4m\5��d��)�d�v�oog�J���{���p��2�'*lV��xM 	���u�Q�:�X�DtM��F�|T�}�B�o4�M��G�q����������nF�������\�`3��Շ����$���;���a��@&�1"����1�_�����4:|�ku9P;�7������g�L�eq_�t6���|O��]�k�}�nt�GA��5"7�1p�%C�߆���a]<L(�kX��T�g����/s��LQ�֫x�үJw����r��.���.T�����U�WU=�
�(��54^�5(�_׋!��"�Is@��Gw[��o�pU����G��ۗ>>�w�'���Z�\�6*��k紉��JU�ԑ�>�:_e�S�T�(�*v3��@���g6lf��_�� ��<��x�
7��m]��Tin�,_n?��Q��M�%�u>W���oj��|�DU�%ߙNI�q�uo�7�'�Wj�ZKh�bT����
�{Z~��u}s]�z�jX��G��U1꾺6�"ዲ������b�>=�$ZH�{$��I2�|����,M{;�����O]Z��V�љ�$7�^���Q���Xєo���(rК[�.`w��Ng�e�C\ty��}g�hq0ď��a��«�����g-��� xVȄ�������.{��V*�],X�0� ��#��r��W�>ejM�ζ�禠]��G��p�Ժ�1)���җ]��zz�>�}�i�#�Q�#�*�É� |.߾�^k���ʹ�
j�uR>MuP댵5��0�s��9o���sѡ�0�68�,(D�u�ǽ��_�I��A� '�J�m���;ܥ����b}���sL�\Q�d��v:��(#���a�=L�y��B]V��2�"��3������&
|&�<��<Qn�� t�8F����3 j_'b*�p�&tz��J��4��d�<�l�8��d9x�yx�h�Y��v����2s''N�l�0o�J�@MeH��.����T�\�/ƸG�͟�����οh���݂>���It��/����P �X�M3����}�(�P��i�
�nY�O�&���@v�L�b�[��i��n�Is�/�)ࣤ���oTJ�4i}����y;/"펀�o�l�12������� ��!ouL�MX�>�&����S]�4���r��
t������Æ�C��t�� q̍�7���N`�ϯ\M������L:�i�_���&M���.�9����~�H(�^��Ϊ�m(�v`��ߚ��	jO.q��l�=dU�u����-9�.V�͔���� ���LYB�
g?�SK�=$9x�
P��%6���6���y҃��v���A��q� E��<4������(�?uP��t�����߉b|*��Xz6����9����|\���P�z�9���St��O
&����+[ن��Ѣn�a�4Qo��+�B�~W��F�l�z\�m���T���[3�)(�P��zi!CEA�6�-Q� CDt+w�٭wJ�e���;<��h^) v˵��MR���7��k�:ӈv��2�ˣ�0&,TAY�X~��`���ŤYEF'~�ͩ�D����Y�;~2hdі-�Bk�d6�zO�]ij�ש��#<�p�GR�(iqOی$J��E��TٹH!^�L��;����ؾ�(���6���*t'	p��<G:�D|�-��n �Wvb풄�3����&U�N~���0��+���0�i=D@���{6lQ���(.����'�#���<!?��%lH���<s��k�d��\�+uhov��E�8�0=�ĥfhf���|SU���ϲ�����?�� P�Ê��Bb���~���Ӎ�-	>���y�l�L��=��b�Ë�Fqv��"�&	�7 ��t_��3�$����̢��T ����X	�s�~���-�L��d0�{��Ѣl�	&���n_/���E�n�D�+<�
���������0r`j������?��0�RwGFms���^EtIM	������P�RV`����8��o�z�Ƣ�ז�=n{.��d���	���<H�M2�4�)�@��+@�������2F�h�d���ygP��	� }��ɰ�x�l_�>���F�`R� ���.�N�*n}��4�c���dG�ѝ�9���>��G��/��H�!찴%��m�j�"Ȧ���������Y�7(N0h*����A_��}{5ب¦1p$��]�ء��:�^�$
/s`{���oC���`ZS�f�գ{��G��Z��k��?���K�ZÐ�!=i�A/����Eu�-"�}�*D��(2� ��Ö�C��Z�F����8�]���#OOx����?p�5��Ljִ�k�+y�9d��W�� �3�X��dw猚ݬ��^��9R<�K�)U�;6�[f����["[�M�-�?��0(�2O�-�.O����_�%s�,D����SŊAM6Z�Y�*�SL&�t���b\�Y;Ѣ�A�P���|��
E�-|����F\�<4��_��\coIAX��^��N)�se��J�t��6�}=|R��dbAΑFN�\�gEu�C���T����A�@Fy�R^s�_��L,]M�����n�]�n�y�o�]^-5�� ր�̩^��:�u�a��Ʋ��-?��
gj��q���RRӒ%�"�%Ձ&���¥KE_F������N� jy�{�$���.#e��$�i� �����ܺ��X��r�H[�f�J�ŋ�$�YE���ڝ�Ux���ξ�����B(kp��(!�,��(��X4}�ȝ��:���ё�-ieMҰ����o�R������b-���@�rT�?=��������)�L���T#}�\7�}K�xmf$�2c���DT�ZPf�ݡ��v|��*�1akk�W�Rqr;�z-�^MՃa��|�å"|aw�KO�tu�E�EtͥO|`q�I��D�ni�$�EW��ș'��v�k���ř����o���K������׫��{��&�T�@5(�>��A!�G�聗L^�]�{ʇ+`�mɳ�V���;е��J+�	����������G����#����� ���侈��;̄&��k*K�M���'�=1�ے��A�'�w��y�:����f���#;'�V��</�)@����dV�TKD���D#񾡖�{ICS-���R�IcPd��u��g�7I��;�gY�c�Ѿ�tt��-�	ҧӠ�,ҧ `f%#Q*@��O��ǫ��;�,�	�\5!2�~P?���T�Ӭ=.I�&�A�l5/��h�t��zg��#��I .��>��:�"�C��CB�|��w6�렢ݯϓ�m�&�4[}J��E+��]�m��`{�'���T0�(c�Е��+őL���eY��sDW�%.��?�|�JX�y�1$N����z
�<�e��d�����{YY��6����D�)s�n\q<W�G��;�l}e���`�A��N��3r˝�fd�Z�@Ya�arP7u:�趜^�ˤ b��?� ;9D��P���d����͓��`�wa2:^ܕ؃R�R�<�h��-�ݠ��������7�S�V��lbP]�Ϊ��TQ˚��43��wX��œLg���g����"0Kb|;��u7^p�<��,a�됈��Xb�Y҆����j�$�����k�����µ�Ζ���	m���([�W�>��a�3Of�Ȳ#��bM$�Ҵq-��5�F��������)]�7 �0<i�IΛ�e��D�������<��w��7�P��|_�Z&���+)@�/C-T��n��z:~(/�&G�\�]:%�<�L\��:B��Kǩ0�x?iI���`�]I�ڐ��ݐ�]pڃ����<�c�\���s�h��q����==��Ov��ɼ<�;�<��ʽk&?4�Yi[�؜�sv��XD���~q.g�/�q!pn0��bgV��,��"�<������`����Z�3�]�ť<�V/iʦI=�f�aLu���O��,#�m�p�dK�I�Ĩ���*�_^��b�n�g���9�H�6�'�g/+��Ej��x�iljznB��Ȕ+h�����M�J�X��fge5pw��ρ����JZ��7��N��L�[�����H
qe'.ج�m�;��7��fQ2������
��?6�x��C*ƷRd��y���kk�gP��֗�U!���R��_,Ȓ�S	���2�Iz����B_�!�xP��y6؈��:.��HQ�rt��ܷlM�W��ѯ]���d?�	G\���l`��V��.N~	��yXwؘz)Ά9�C����'�
���?��}�O���~����P�޽�H���u����|��ր-g�6�k�Ρ�㖊9�څ��yXU�|����2��q\�̜�ԍ�"��Ֆ���i�K)���%qk�/��]\t��aq�~�q�{ȓ8=���(�o|míC,���N:'�˅7�xF�JB'@a�A�E��l�����76��UN���%^W�S�Ij�������xO�.&..v
� ��^:z�Ig�!�>ɲ�}��K�"���*�w ���+���D���n�RQ)㐼ދ�X��U�6Y�.EQ��UR�����	�Uv��\i���[%�5})�>=�gP�' ��� ��nU��d(�EL�
�N�Gz���U���jMy�[��"n�l�RS����3Z�v��~���R�4���wo�r�������OβHR�1�1.��ͳ�c���O%}���@���%�E���2�"�Aݼ���h R��AB�l)~���a% B1Y��z����������u=הF��?r�@�򹲏��d�̧�#�з����|�R��Ҕ �-�A�]xLM{@[tZ%!���il*��S�%��Z�E���ؾw�JW��Wu��h��7'�B���:�z^����	�P�~���|r@O��0�ܩ]���D�W�����Y�r&X�_9����<�p:�����?WԮ5�y֨e�C0_U]ȡ��Pټ�A��������'���rG� J����@�T���؀�K���%!{.�Uֽ��<�M��}g��0�2zk�D��H���]�0�'v.�i�#��L<�oH�e>���RBHl�G��ޟ�6���gx{�Cf��O�g���BrDՔ�畑S�1�y�����*���@{B�`���n�X�F�_'���^�yp��Qm��%���\��=�q���8c�芮��wf����{��WE�g�����K_��s��)�*|�Zƾe|7;�A����p� ��v�=�\�.�I�~Y�e)Y�vt,ɋ���yUжx�!u�[K�o!^�y�$��wzK>(X<��C��}��~�v>�ɕ���������J%�S��5]��p��	BX�K�d��!�Y�.]`��|��E�y�m*�v��F��������d�� ������G�c���n�$�[3\mI����a\���G������� X�"K[ݩK$s v�>
���X|�])�S`�ea!��.�f�@a��@��)N	���i���[Ӄ�_���+_Za+\��	l�5Q���/oc�|��f�ܯu����@q�å)K4Ij��W8 �b�9)NÞ$�4��->��V�20�1�lL�h'J�?f�������X0�3�E�J���wp�4�ˁ����SS�l�rfȲ�����3�\5�/�yg�w�X8�W�)2^����-�A_P�#�<�%��D]fq�td��&���lGۉ ���땷�3���+����������Z ��}��1���}џ����(����
n]����7�����?��Ո鍳"tF���E���5z�C��{_M|�	I%bQC@��4�i�F���6g���6t�j����(���x �x��R��F+�>������m����6ݴ��N@�	W�� y`��@�z�ZI:�	˯��L�P3�J�W91Ҽ�3�,��Ul�'v����lW��I)l�Ķ�g�%�� O#�X:���܏w7R���i�y̾�	`�*�d>[xۨ��O��^������k�#K����_&����&�m�$��3褩��Yb t1PG�_`��K�w X��j�ڒCFʍW�ь��U�H�ǥ��3㜚��?���n`�����8��f�Q9������*����e�E���o�/��-L��M�3���q!s '(�+S�w��'�+�U�
uY჎%�t�
A��x�>�U$:G��S-��i����g�0��5��8��Eǽ>�r�q8��g����pE3���젟�*�������f��7�5-�Uڎ�\�3~��n�Iɠħ����kX�e�<Q�Z���@#�(���Z{X��,�By��NX](��q�]o'�!n���@?_�)�����́�"Z���p�� M#�³SL�U�0.�����O���ϥ�jĺT����+�s��<0v0��[G�Y	�qS�b�o�]���x�3Ư�TY}��>?�{�+��;g5�S��m�n5�x��o{"F����dN�+ܖ$�^^��Y�3x��!t	�=��Zt_A��׌[�䋨�.Z$��E����9P�"��.XX��������,+�'=_殃��1�,����ʿ(�.�4����ݝ.,���]�!ҩ �4�Kw��t�H7HJ7���W�_����n�s�ܹW���"tE�P�R�&9�JY���������w�;�d����)��7�r��^6�;��8�X6M0N��*�%*�+}�~W�/�d�Q5qmG"��%���^]�� lJ�cS钙����!'y��O�׵�e��H0h&+"W�1�P�@�?D}8e:��X&	���J�|��3%s���nk�}xv>�A���?r`�0Mp�+w�(�ZF�ǘ���/��u�k��;���5Jy�(�
h�͍gN.�3��o�uI�+��uut�ɫ�:#�DMC�U�:dnǾd�6��ۦY�MMR+�L5֓�)�����S�__i��?��?�c��O���NJTO6<�8���H�#����>��$�=
�h�YQ�K����ΌƇve&?7�6d4��z~� �.xh�mb�ޭ������݉~~e�被h�_�J��Y��R���᧳�驀տ̃�2ҝ���#���Oys�<�&M)�� b
+��K�G��Y&Hǎ�Ȅ�)m"-)��y6�Uj�x[�Z�4��hp#X���	���!����yu�P�m,:��Z�)��	�Vׁ*MoI6���W[%~k���#jē��S~� ʳ����'~�F�&yK���Y~gi�V��V���hb��;��.6�_�ս�Q>)l<xr9URbࣛ��rlJ���O�G�:��{��}�����mU� *�����}u���VI���PM/t=���9�F��ꬬ�VAS�|#�ݘ�Rm����F�����N�b����%�^���K��F�����b-K,3�����.���C�[�do(��28@�#��bQ��"e���j�Xė5s̵�Ŵ#j�)��*a|Ո��ѩ.��vx&�h�v	P �w�W��Q���V��MŰe)K�����cO �B�O ��o>a�t�>���W�W"e�<LJ���a�����{�7�9b���z�PJ�w*s�#D�?�X�~���L��.z)m��a����{��|�W�|�zߐɼ�6����+Ȫc�!o��G��$�vU]�������`�FW]��W�~��1֪y�96m��hm�������9�\=�^��Y� ��ܿ>5���S��:���Y������[�Z-WE�?�	�K� ���)m��;q
�a��J�Z�ي�5(Es$)����<���PKęn\e�{�����q��Z�����RF]��"��ac���((�B��g�|p�&[���x���դ[Z�{a�AdÕ�L�x���Bh�%k��~�F����P�O��	L&ΠQ")}!�	�J,||Wnۢ��B1��6|N�]�TJ+��Tu����n����	B�U��.J���Wjɫb3C��ѐ�,Wq�z֕y�A�����w���BѨT-�=+	]Q\��=i<y�\�k�e9L&�����kq������)L��-aKwD(��7�?���R9A\=յ��m����zЯ�T�-+5 ��yе��^]�s	�џާ<�(��T��\;XǠ�<�����0�4�"Nd�p�صa1q]W3Ol�����~��1��Ͳ����_nv�_	���.�[x����@���N��l�$�����M%!�li�����?�0����L�׏��7�$����D�>��>#j}3n��f(J%�c��2$)hDD�'���Fk,��YW�!�1�.���mƙa:g��OV��_I(�����\�3<���X^��-y�c9O7���Zl�J�ڍ�5��v�_��m�A.Js�5d\41�à�p��+�e=}��ȑ��aX1��2��uY�OUi�Ǭu��m����FD��^������v),���Z8�Ԉ�.ll~��H�Lr2$��/0%��?!���]16E ������g�D�w�Q\Ā��Y.w�X3�g���p���ۛͮ@�i9�2�������C3���`x߶Zjv�-ְ֏t�{C�ggsR�x����f�g��b~�G�R2�oM�:��๋����!��Haɧ��ߨ�m�����
pH�=�y��0 �e5�8bn9[g笴� 2 �S2	�;r�`hX1�ܪ�0��x�z�_Q
8��&.5MO�ǥL[�����c-]H�i�ˑk�g*�M��趬�/�)��&�4m#�/��ƍ�>����m��=���QG�#�iY��DM�/hJ'�9�b��E_?()��~��,"��Mh���E��<���@�7��#S��+Ze�,��D���I�ql��/��5�޲�8�p�}��0˃^�������5�c����(P>xKwO��Vl~|<I<6u�e+@QgzjBι��u�Q:�E8k�ӈ�#w���=�%�#pT��e�Du����^_qp�s1k��-[�S�^8)M	�$��w���rÇ�ؘ��"���p"&5<���-Z^,����ף�æL��$K
�)~y�On�8�~i�4��ݲQ��o@�ݽ/l�('�ia��]�6�I��=m���FEC�F*z�2'��aR�*��G�l��r�5�n�
u=�э�y����F^ �p��yRV����aJ��	�%�c���rb�_�җ���t$����$���>y�V� �8���G�e�`��w�C�Oe3�#]�Ǻ�+������(��,�jʷ�iX��:b��9\��I�]7Y�˹��pe��bLc���vT}MN��ȅf1^�"=������!1��ۂco��4 !R�6rDw����hR�'���̞>�E����粃5��ݐ���ql@�`'�����y�As��?/d�\�?(e�n{��h�o�px�v�t�;�R�	����J�-_y�d�lZ���[	�6<��Vi��f��	@��kO��,	JSdޣR<��ؿYDB��$v%�^�o�kx�>:��Ρ�hb�d}el@���
{c5� ��@pR��%{�Y���	r���}J��_�[������$L���":�lx����AX.(0Kq��']S%U�_g7��`޿����f�M����?]<?��صe�ꨃ��Ig��/�M�nU���(=S���)/�����%y(CuMnH,TlaB�Xч��'L�%�>U���������ѧ9�)�o��SW�Y0��\��F^��S��{l�����R��a%s��3���X��w\O|�[^�f�3�}D�:���X;������AS+���z��C�?�o�P�>��X�W�8�a���A!L+���/d��\�>��RP����B'7�Eg��O���@�u_�|���C�+���s���ד�1v	�����,�G�Dt�h�+���x�8˝ZF�5���r���s>e�t`�;3����Pӻ*F���;O����#���������J��H{�:�X��abʣN� ��2<����0�`~�W�?<(����M�"h�*ܧx`�B,\�2���mr��W�
�!��Pif��4��<��y�(��GY��E<�3&�#Wm���;h����j�38�q���a~���
�a5���,�֓�y�V���r�Ƞ�cK�A�=Q�T��)�X^��}�߬���$O���z|$�PR,Zz��Do,��GŻȫ[�-�4�/|hwI�u�F{@�	
�L�t|�-p���B� R��W�Š� %��@Y�V�Y�ϛT˟��߇���*�n�Ly�V�P�k�LG��V�J��ǻ�s�_����Ɋ&��y5u���N1gI��ϳ��( /�u�&,�洭N��۰�s�˿��pF��!7��{��~���{���z�~�_:�<�z��uL� lA ��d����^jtz���F����7xl����!&��7� Ҳ����(���6/�=m�O�'*1�!�c��	R[w�Ǎ^��x�[�%�X��r�Rzk���`E���M� �/�Q^��e��U4(��h���<���L�0��b�����"���k�!��ݵ�#�R��+��f�>�PU
�fqVd��	�� r��i����J�eU�|�EL����e�P�g^TW,�F����W��v@Xg_R^�7�Y%qvd6��������2�(����gΠ)���u6�½�քܓ�'T�I]H��}s��+u���0���~06�(��}�?�H]��1�ށ>�f��2�����ҿ�($�T���U���v91�{��yz�����qt�HZ'-Q����xf�!��u�.h0��m+x4��Y�U�9��;��
�2j�����/�����R �b���N��chO�^t�X��s�ʏS�l��mu��dZW�F/�S�O.b��vB2�)��	���eЙI��<`:~(?���/9��3|�Y�p�'�D����&XFA�z���Z>��)�>��]�'�|�a�u|m��WB7������j<�<�ru�EݮE�m���n4��.n���0��`���tZ���I�3"�T2����5�.r|��1:k9�6��+���V�!����	G���|D������w��B�M}j��X�@3�A~�p��I��R@K�Uu�+Q��ĪV��y�VF����Bh�X����)��{�\�Y�e�S���6>��2l�JPxt)D��|k���(=�x�>֩��4je�;��3h���5�i��N������r3�b���?��f���Y���� 3('��A}h����^���Yn�5i��N�h\��$Z;F|c^�b�B����TW5wͯ����"��]�?�!j/v�56D�}�Wz}�5��!��G&I6�EޛVH����f`TrHU�UK��ш�oЀˁY�ٜ-�>��gj.M�bk�сU-Ƃ�
��舺f�\�ݼ �����B�=��'(�Ɗ͞9*.<�'�>KPSѐ��%{9� ׬��
d+V����;�\�dEC�i*���i��ПY���@�/��7��4���M@U�V��Jg�I̎��o]�5�)�/��g�܈o6ˣ���� 2ȳ����W��'�����'��4_���~0�ۯZ'1O�2mX��;8�W��(~��.���)kN�_�q�8��L�nQ�Y��ME]�+��z�c����W��2v5M���ͭ����+���E^]�=e|ZC{޷S�l�1��_1��}�ڔ	 ��O�%X'd|������1�����sꐟ�
����?�lN���Um {*�L\��9+I}J�1��"�/>�v(�qz�)e4(
�~�~�-�q���y�Fj�j��.������d��C�s�"y�=9�a��}�X�Ļ��G�{�R7���AL��Q�U~���/�ܰ'(-�f6�T8�)��댣�e�k�Y_�ǧ_wh&h����x%
�H��æJ@_zT�>v��߷��vg�}L1P����U�֑{��@��F]^��������Ve�4j�D˾�/C�C�Rz2Y��4��x���[�d��!�|~u���#�C+�*���n!����ن�]�D;��6`�CܮZg�m�;���$����j�{����#Ư��+�����H��x �A�z5����E���b$Ó�5~�D,�y�T�ު��`�����.Z�Қ{��ur��N���)xk0�G̽h����V��m;�`�@��,�s_A���k�QQ���)hd�K�86�@����̛��80��z>�'mN1+��*��������Dٓ�`,��zLTc�O�u`�-)�`��;UW�U@*�}��-'����\�\���$�j|j�<����ʰM/n�6������N�*��z+��q�Np��sӯ 6�yĕ/]�-^�N&ƒ������܇�Z��j+K��A�[#gP��^���`<q�)�i�=�<�|�����s�zjGNG�x�2G�kV���Յ�͌�9�p�"-H"��n��[�]Mn��`Iy���!�=�O���!R9d�]΃s� ����t�����[�N)c<�I)���:$�X�k`q�x�};�1j�`@5�E���yƽ./)p-Z��W��,<9��}�����\�<t���G���f���&�Ժ��U)U�n�v2�4k�
�9����t���WW������!#M���u�n*-��o���*+(~������:՞9F5p��c�1�.�N��~z�	��ڲV]/%�b��{�Dz��l"n]E���1��/�SOj�rG;�>fd�\e�g��p5�����U?�(��仈 ^ ���A�5 ��X�1q�kHEX��`�5 F���4���3�r;G�1i���vH����7'������g�\r��*B�%�)�#�m�����>�l_�S�k~RƦko�}��j�r��P�;��w�.-��-��f/Btŕ���H����J-l�'V�GΥAmEc1�v�ɲ��Ȇ@�9B3�K���?�m�������G��Jp����{�T퓁G�-1�R�z@�Y�}�t����u�����.���E��aL�r��p;��y�6��bH'ɪ�.WiH�/��p��u��r̴�����>jy�n���`KU1F'|l�ޤ�^@ֿ{�Q�24v�L�qT�E(+>��8;�����'��	��	�T��*r�G�\ݬ|��3�x�	L߆AV�+��T��a�p��^AHW�
�H�x���|�ƞ�K�j����%���*@wqm'���_-�۠�g���*������J1�b2VL��`�V�����\SM݈e}���ļ�.�{R15����?�9h���ᥥ�c�y�N���"w,8�#YYM�ɰT�KE�i�o��I��]_����U��+���犠9�!�.�%�
4�W
t����Rz�j���Xi�!�@��T��\��!Y#�v@	į�|�Ɩ}�`/8�?�#�E@r��tvk���_��ˇڥ�)��`>� 7��r�Υ4�����c5;�(��~�4�{]9>��|��AM��P�'s�d���Ċvp�T�����!�<�P�3?x��Dkp\���'��/(*X:<d�P�?V�ӽ1XQ��L	��4�0`�ڂe�'�(q�	�� �}�'��yw�h!�#0�,�4��V��ኊ�O�{�q�g�5�7���{�iOa�`�t�@� �f�����7FZ��iL����9S�@*L�k.����0|4�4'L�~c��h�o���݋�9��a�������ZZ������p��ȥ��H���ׄaGELh�@�쐋9�ҟ�[���V��Zo�s7;��7uZ���P���Sb
��G��K�m��?d�$5&�؀S�.��8$����JF����p����Dl��5������r����+�3C�9Y�\����κP��/�kG����#ݩ;�Qsʐ�J���G���^7iN1��n��[[��T*�W��S�h�@�Vo�C9��-���zd�-)wt��}'��"��tO(ɝ�+-�
��3V~R��+���R\�br4??�Q�<���}*���I��"������'��߳V��}��j����`u~�T!i��N��莪��P�|����\ 
���cy�^uIh\����!������f.[�dV0Oܘ�+F<`�G��f���~IE9�j�n^kD9x���^A�<�H�Zw�T�H(���E�����?.�8ے�e�n��I����� z$�[�l��xUn�ʛK��(qDF�W9L���'�>������2Jh��{�����ᒄ�)�A�Xu��g�yNKnCa�@�VjKJ<���Z���ϗ���d���K�:���U���f�b{����}Y�Y����[E o+�%�w���*HP��%(��ה��nla�^_��m'4Ut���`6��Ef��j`�H���ܦ F���>Cs��5���ry�s�<Cr}"׳�R�C�4�� �v!������v��(\+�)�Ю1]��扤��"n:��ő��%������ ы�ߌ���0��,VAga߽��@�q����f�\����������ׄ�X���RLq���/�ښ�����W�'���4�^�i�Gd��K_�� p�c��C\6"�(����7Q?��,�Q"i�����[�t0��1�g�1*�5 a��������S��[�E��!)���5��Sj���ЖA�0���^����P��V����̻�J�r�7|�|���]\�棘1�PV"NgV�� �\MA-�3O������a���#��$����k��)�sN`G��>]�[Ŋ������Gg�Ҽ�Q�ì)m��?��,EH�)Ŀ�8���k.Uu��T,�D�L�<��3�+i��R�V�sK�R����������N�U_�,H�/jO��0�A�w>��Y�o�s/�*�cE�Wb�Ko�{��f���-�j�4w��o4�eA!�%b�A�NghW����J攴�I� di2�̯g�r�bs��A�%+�D'�7�Y� ��<-�-���7G�������)�U����B�7؎�UWZ`���Ґ��$�j�?+��H鐵���,FTK3��^4�U4WKc�|�H���T��-�fѺť�������.��������q":�
4g4BP���o������_�[?�p>cGM�_�!t5w)$�v9
�C�2��lԊ��}�{�!���>�����/KjOa�4t6�;%F��\�ܬSA���6!�ڴ������2�SaB�\q�Eˎ_�-g��_d��ŀ}�/�kj���C���C�m��tJ<��c���,���~�����U\�+�)�橚$Bm+��C�?v�>)T�
�F��^:I�
�W����i�>�������_$t��f���[Ka�%���n��|��i�P�[�g"	Ӭ̑��ϙ���$:o�׸J=g��F���Vl�<�=���0��]պ�����j�S��M�1��ʟ��7��}�h ͹qy�4�'۰R�=eu1��)��z ��[�'N��
�e�j�ߜ���{J[��N�P�N|�d�]C8��U�͘� ��;_�g��L��o�%���F�������TCb���h�P"�^���"���G	1cGSEѸ������8j:���\��Y����	]ĉ�:b�r��w��#�I�^]Mv�NU�-h���g�1�ER`$P�I^���ɕn@�5��$z2.�//A�5��R}-����O��W���d�WeMSTkB���a�N=�xX��.�9��z����c H�f�B*��p<�[Z&�y�;�l�sx�YK�����r����I��1���h,�%mx1�`����zQC��Ű��s������`�AYt�Q�тJ���X�ҡGd<9����v���@��((�A�Y����Ka��jѿwaEJ���,���4+�<�]猪HxRO��i��3
�J$5�ׁ�vGot�*ͮ�g0B4;P���C*d��F��'�ajg
vsyxʂ�jp����>^�����UO�)��Ldƫ�F� 5��ݡ|��H��CU�«�4.�bAs&E�	�z��"���ۙ�1�`"�VѲ;-��<�ˁʛa&��]��aթݺo�>���wB��F�d�+,�`�k,���c���ַ�G(�l{�G�x��]Њ[UQ��T�-0|u��J���;���5R���o���ƴliK������g1okh�Wr}p�`�,�l+-��΃�u���fˡ�T��h�|�$bkM����L`@��yu�>��
o<��7K(F}�R�;��K��¬,�/VQ7"i?|�e�5t�\��\�@Q���Z��F�<�Mr/hX��fTe�� M��W�*�l�I�#�V�@rΧ����ﴤ���n�c���J��P?�ʭR{5<��8��QF�M�N�X��d��M���1��:0�ǫ�ZM���
���́4�N�m���jc�O,�2'�(�~/���`����yXc�!�~��Y�p �p��[v�F�קd�҆�=�W�i�:/�����
�Ž����=���j뤹'��~.J�t������zhxJ��|N6��?���v��G�G8<4�r!�ru�� �������i�]�>g�}x��=��t5��̙ftAf�4ChsN�id~����������:�����5��M��l�|�.z�O �O#��(�|4Ъ��.G0�d��ß�&a�ȣ=�
 �-�x�[)ѿ���j猛$����LSR���@d�œlc:����y��gYW����QG.㍠�X?;[VK�wE�#���'?埕�$˖�5�QX7/���C�?�ο�&����,$���K_{�mXg�w�2[��(���RN|����҂�����j��6V����4N_��n���S�R�*��W(���媩�U�]?y�bl,�ٔM����{9�.,kZ���sė�²e�/��%)%�55Ԝc'�%���hR�pE7�N��ʄ)�u����� �W�m�����dPq��'J�]�Ҏ݀T��gg��R�or�C�]fKw�9�#C��S�_*�f������g��I-�q�-��F�H?���vB��� ����Ջ��OuCn��F̂�����Zpш�s�����
��67��x7�k�n�D���s(�:��<Ѩ�p�'����b�B�*6�2����ʀ5..����7J^��7��Ǒ9ȹ�e�3�x�gODҾ��ȴD�h��;T����c��sf�A���:B���c�zG�5�3�-�eq�I=����Y�i�̉YJi��qImibN���o����=��}횗����e��ܽ}Z��&:9��9-V����},���bDR�I�]f�C#Q/�q=���T�U�uu{�݄9gA,�qP%&l�ڞ$e��a�`�M�����<�_�q�TD)��v|c�:����O���k�&��������v���5��� ��igG���\R�H��J�2\z�}�B,��~�>�6fz͗>�l����������|Gn�m[��ΰ�~�+bR�a0W'�(멳p����d��'��u^���䬂r��(����?��>����$�(��t�휉-��fRf��d�YhX$��uH
��vMPJ��	�d{GN�Ej�4�=7aS���������OR02K���J=y�b��p-�*�H�o��ki���c�L��D����i<�0|v�xn�_�M�o��TuFx=�N\���a�݀'��ҽ�6{���Rڤh�-���9�6/��K{Z�{�!�B)sX�_�'���Ì����S�˭����o%GG���Ӽ`ş�M�����c�b�e��<�%�<�\``J���/��B%{��m/�2�]�׮H�l {����^��_�aݱ��)˷σ�	�Ja�ď��BG�c���6>RL:�v�L5E�/�(��=ha���(�����#���7�Գe���JA����I�GSè5�5xث�د>'�T���8���s��k��	�����@�J��2J�@?T��~)�+R	��y-u<����{��BN+�Ş��g _��l!�txT��>�������5��F^�2ko��iǴ�Ga_C~��[M����rPGXs-n� jQ7dQ��ǴU�
��z-�f�߾�Q�m�w�&�`�9��K�˗!$UD�ܓF��d������y���*p��h����j����,�W��C)�+�wO�&o�$ڱ.�Of�`h?�r�ȧ��!M?=@+M5ĺ������=>�Y���M��r�)
yD�bu~�Ѭ$0�����J����fhޓYT!�juDii��'� �Ƃ/��O;s��4Z4����2�Q��Wqh��@���f�Fd����l��s2z)<APz�S���-$��a�� �Ō�TBJ��'������
da��ŏN�L�i��`��V���0��a�*#;�*������|����B���옕�2����i.XNN=��5=�ܮ��T����$*�B�<Q�@ ծ�?�}Ki';�K���!!��	E3b���'~v����ξ$5Gd�a�����e��͈����~��lp�޲�����tG�����	�uT1��P6d��{�Z*�A������Y�@sqSN,���񖺑	�/ M��o��y�ݘ�����B�>Fꬬ̻ʲ�9?쥵�W
�Q�d��/�$�˃��U�8Ija%߽�� �믧��C��f���$�V�,���:��Z;�� ��H����GP�.9��I�51�ƈ���LW�R!`7ٻ��5V`�`3쎊��/����Ω�L+�b���NYM�$����� uXn�����Q��吇A�pM�ENR������b��p6_�\�/'�,?Ef4"H�PRHS�T�����X$�V�J���ࡡ�{
��z4ti5��8��U���W����u�x<�ǯn�@E�A-Os�(�+=�!JE�&~x��=5	�2�16G\iwNN�DE���S,��dᩗm�NP2T�9T7d��鱶N[VkVw�������M�V�c�M=��ֈ�M�@o�T5�;q�wj>�Ն{a�H5�C��{�����`��sc�J]�-aI[��o� W�8?��|�ۻb�d�R�X�!$uu��̮��㱑

�
����8QL,� ��"���[����4�5ZV�<<ߥ����)�6��U܌s������\��f#��@Ts�
d���8���):	@m�{	jYȃ�;]���Vd�rR�1g�z�|CU��Pt޶)���l׷/'�U���1�>h,�����Y�t�/����7%�H��I�&JS��X� s�9}`��Ky9����t����S�xj�Wv0/w�r��T1�: �X�������&X.��<��(����L�� �>���Vֈ��hU�/�6��Dk(ܮH��u`H��&���2aMz�8�nJ�A.�rU�N��FDB��l���4�KJJ/�;���\0���#�U��I�S���Ql��Z�eW.<B�.O ��^�c+�a���ZC_6����꫖�j�Q.#�.;θ�uoIaA	�'�[���C��;.+vR���P�6؄R	X:23��L>.hT���s
�JP�� q|b����/ᛟ���$}sun���p"��*�W�Y^�-��7O��
^�+עn����m[r�i8�K^r��q=�P*g��B!��3��Y�=�{wkU�4�1@ׁ�8��jj	[7�R�A�W�[�g0��٦z�^ y�C'�(�-ѓ��cM3�}�	������p��K�v_=�=c�J�_1A}�CY�P;�2�)OF@�y �=s�0q1zT^����~�G�p�nS-'?�1(}�(��N=[s;�4}�С*M~���P>�:��jP��N����Tl�'�E�Amp����z�r'rh�ۭac��@����ܔ=w)���v�?��)|�+�h)7��Y���ˎ1�<�A�`����&��Ǘo{jھ�lT����%z���ƭ�[ ߘ��`��B�&�Ĵ��j��C���ꚐT�W:��EѪ��5��+$��҆�&�`������l!Do��J!�=r�d976��YlB�$�V�»��	
�*n�D�Sqz[�sf����ֶB�S&��j��}MDM���Fd��s"ζp2'A������B����|�[_��(sjj��!r�p:���Ü�ssF M����Ylc]�����Xz�=��e�k���� x��a�1Z�o����C뵳I�3���UyX��+���D��.��L�l�u�B�c]��14m�*���aZyt�Z ���CxL�-�O+��fg�Tc9�X-8��r4a�%�|op�%c9� �ӊ�>��ÒFn�u��bl �����S�ΣJ��zU�o�w�1�ːs̈`qh�)
j�]�ةP7�Nu5m~|�7T)Q���Q���ǌm-m-W���r�WZ������Ssq��J�h}&�˘,���3�k���-ۉ�Y�^c�|�b�_k��.qb�6��da��oJ��������вt>�
��$��ۥtQ�N]�Y9hcWaK�MPу�OH�[���1��3����'��$�X{�O+�n��ȭ�טs5r(�]S�����XM���Q�j�)qu|�c����� �{���ǐ���U6EJJ�>��m^u��w�h1������'�ssŞ��8Nl����!��0�LnV���.�g��p�<�U=�Q�(���L��t�ԗ��	��ػ�,�6�&>^�$D�$C�B{\c\臯)7J�Q�����cJ�*	5㥤F���B=��,��hB�bd=�d1�1���R�*�(��V��� �S�)NFs=-j8�&�+]h��4y����>�+��F��#�?���y*�v�.k���	��=�dS�W���繾�`�2�^��@�,� �o�]M4���C}$}c�U��eH{�ʌ�����B�S�/�[;Ӝ�)�0�(@6wb�rN{���g3�)Xd�wk~��ܮ3TQI(*�*I����ȰH�)�mK1kv«xL�t�i��v��M��P�zF\I'vz�h.��Jv�n�ݷ-�����?ە�fq�[\AKfc���`�'B�V�;��R.�1b姊R�'��֊����p�9e��85�Ǧ
�Z����;�>���/ �����hZ%bѯz���~͑<��Yl�v��f#��	�YOU���0̙�_�^��]�NZ��4ZC��f/A������� 	#ץtB��t���zg�y��(xH�z�'����c�/�4��4?w&W�UV�q���:E�J�u9���ΏƖ�״�ccu<U��<i;����0�A*S;���/ ^�,�d����������U	�g��l�M��g��.�xu��o=K�+�7�����󂚡���ܹy1��F�.("l��? Z�Z�cl4���H@aN���ȥe_�����x=/	����/J$5�-������q�K������I$���wt>[v-����,Q���݅�]��jL��X��_�����(e�F:�ڄaƜÉ\�+����05g0K:=�q �\O`oW�h�D<�����f�$�^�8�K��
m��{�y-bNY����(�Z��6�����b9]��.�e:�2�z��}{��>Q5=%��_��W!ZV:Ȗ\�ޜG%�d<�>]����� �7�¿�?��р�D�Z�"�Y܂P֓ҿ\�k[���aPj�y������Ff���{����O��=��.�ٌ���Sձj��+�H޷2��������~z����DKڸH�J��|L�/��Z[Oˢ�
q�xã������~,�� M������s<�Ԕ@f�x�<e����a�_MS�#��Pԥ���ޞ��'*��qj��ҕ�M�^t���I��'e�o�mr(�r2S��^<:׍j�u��U)�)>�����XTʷ�b"���э���7�R�O�9*[=��ն����2�'�y	[6�J�i1��	-e)�Լ zoW� Z<�*-�͙�$
����IH�PK��K%�֜�Im���.~K��N��v�����0䌓*O�m�̤�g�J�U���k�=�@�|^��:7Q?������+�t)Ϣə됚�}��BP1����)�I���1�G�ǃ����IZ��{�R��%·�Q3j�[Az���N�kc���9K9T�l�!����NA��0�˹ܩ��9��{��� ��d���6��@�{�^�W̯���Ą��>�e���){�h�\�~~�{��4���Om756�@pU7�N���ͥ �w���v���k�_�E��89���ha|P�C�"���	�_Ѧ��������.��$��|T��V3�u�zO-�6��[����c(Y!c.��$�f	sSxx�jk�UҙEX<u�p;x�ӯ�.�L��]D( 5z��7[{_��(��ä��ut��Z�G������؃Zg��7�m7cNDԦ�4�Zy�Պ�5�wG� /k��~�K�C�H}�(ɔ�c�Q$4,Hi�|f�J���1s��I���׀AOab����ILA1���47�wǈ� �:s��E�8@�tA���(�����"N5K���F����Ͻ�gc�/��� ����Kr�.7P���}H(�0԰��"���$��[�m��A��!"�Po^{j~��ǵ��1Nf���D��t�HҤ-��"����o�{S]RY	e�t8��3��)���lI�'U�i^���k�>�>��W�Y����FJOFgv>K��߭rl��{%WEa�t�VH�Ƨ�M�`��}���I@\��*��F(�/��W�ʩ5�/ ��W�yv:��uɌour	����!��.+�l�Wpo�t9w���`�JC������;˭8��]7�.�!Hpw����[�Kp���ݽqw'w�{pi,�7_����[cT�Z��\��%Od1�`岺Q��o#��(�*�	�	=dgCt�� � aF?Z��գ�E	K��C��k���9�s��$[��X�m�z,���|�7�7�D0��$���T<�&}�1��\�:zT���3�����i�����qw/� x���o��(毢��d�(s� �+�)��-�cJ6��b��N7ZDF��V�S,��*�>;A\tںU��6�*{��H	�j��a_ﺜ�s*7�y�*-�l�[G(M�1$O�1��Ĺ�e��n�"#�ݜ���(�m���Μ�ވh������/?N	�I�M�Daݷ�(t���i�T��6�$���V3��?aw�^����h@9_�nN5��ڧ�%9E����J�oNoy�'�����[�3=�A|0kډJ �i`Z��7��4��ޛ���	J�I��s)�شJ��_C<>J�A���+&�[{.�4��9����~��"I�^:�=��|H���l�Hf��,-�V��c��@L_0`r������D8~`S��mi�N��֐FN6�ƶꌘ��D?j�ze�%��h��ب�v�wvh��TR��V����� ���J��;�*��B��4���9`����0���S��}x��ZU-�r��fތ���>��1���T�79�2��|r5�6<LZ���Kݚ�%&hT�Cуk!��S"�]��,H'N$�숋r����KQI���ߺ����3�Z�m��M_�pU9T"9x,�
1|'�%�b�:0�ĩV�:Vpy��~C ������~�n����ZvB��pP�o)�T:�5��Ҫ���z�oN�.n�$ϋ
�<]pN���D���&���^��9��Jz?	��g��[�?�.��$�?��=;�����RE�������=��,^4Y�����U��� �}v{���y����ċ�պ���"yѧp�k�/���d��?	0�x}�4�i�8u�װ������Z~q|���X%���[�R�h���.��;G��r~[����&�"ф.;���~�/��sCMؖ�<1�����Di�Z�"zl�̂�����Q Y��²�z+����G�ݚR�UQ<uu��@G{�����#��5�9"�]2��r�_����(����9�}l�����lsR�y����p���D���rHsG��d�\��E �(�L��DYx+n��eD�M���y�4"L�J��|'c ��Fe�k`2*�xJ�2X[�O�\��+!���rv�d� }�6��[�p2P]>X��P4���7��������)H=����H��'�k�@k3���O���r�_Pc�2��r��U(۪)O*c�[����m�eQ?�#j}:���7?�9�X\`T�R&����Q�����L��Q�o��k���41w�>a!�۶S)�Ua�r��
q�ƪTo�}]�3���u�� ��{�E%ͦ��lT�VI�i�F�.iG�5�:L}�u^3DH6�~�r{Μry+?�X���Q`=7,ʶ.O}�=���d<9xzz�ZV� ��۠�%��-an@�w��yQ��\*N+߹���7�ѷ}p
6�ި�{c3��)j��s8�0j}���-J�d�D�a����VN��������T�R�T���Ȧ��
?O}p�ӓ�2�˒b��/�N!�VH$D�P��J�/ں\�{�[ky�߆��@׶Bܔ�V�3�ĨT2�H�yOyzf��t~�F�W��d��s�c)��7��؅c��6?R
�����Og����q�n\q��,�f��J{�)�ې8z9��}7/vJ�`C$�qj'�m]���o[�"�GO��>N>��s[A)厶7{�z���ϖ��?�?�)���G[���ܵ��>\�u96$�����ؾ����Ƙ[�ǯ*7�{²�x�;}>X�t��4�ZB�t&[	H�� ���E�c3+�Jmm�#���Qᎌ1�7{B���'�Up�|:�.u�ew�l��^k+��v˙#h���H[vV�;��mf��P�����4�C�P����0��$��؜�IB�ۑ��?�F�Xޱ�D��-�y+�KקX�W@����b�x��ekLw�c8�����%6�%^|�72@K��Tօ��,ؚ���Ӿ?r�#��+J�٥<P�<vZ������)�YÁ���0���WE�\�|C!�S%��S��B\Szڈv6c����_����0���32�������٥����Al��5[��sV�������Kw邾fL�2��裑��e���v�:��tj:t���
\K�[/2���\�^S�w Դ&ށ?��q���[,<R�M���.��~U���s]ɉ�'A�Yq&�f��j���~����Q�9=�&�,��ߖ�Δ���8�Ԙ��ʹ���ñϲ��K}T�t�V���m����Qa��X��Կ{k�!SL�R������>�9�{?���w�$qzH��v�`�T�N�G	�Q�����w�23{��ғ'(�����)�pEN�D�nXl`�qF7����g��	�p*��;�â]L��m~�>���I�q.����I����������*�<�������t.��%�6���X�n�6O��].���CّH�*��'Y@��?;���{��$l�Y�2��q�|ͺ]O�@wmn��mJotS�h
,�g��Ǜ�A*L�^��>S�<���?�d�����v��M��]�ν�Ei#�?@#�Q�3B�l@v�������KK��CY?�K��F����EB���r`K3�woh_+A4')�v�i����Q��F9\�<]hf#��I�͒6ߥ�<�8������u�#�)k�%�:��ג��p�yR�E)��_g�Ue�nxr&���m��RU�,�Ph�x���$�#�~L��Ly ���[��3q�9Ѷ�з<�HB=U,Ѡ���(L2!�.,��$��V�x��ʎo����B?�/2��)���^v��.�K�A�,�4䶙! ����^[�a��"^㇋3p'y��|k���O(�~��I���>?$�\B�J�	�+u6����������,B���-���h	��g�:˅�c}�q$��	�eW~G���x�n򓘵)�I2��1>E����eE4���ΡI+ ?�'�~l�]�/�6�1�	�LQ�3
�r,�����[c�&�Y��0V�1��l�z�	��~yyE���1k2��ݍ��0u�-u���E��𱻦�-�#�}FICd�c�2s���� /��Qˀ�K�ѣ$��d�9͆ f�lj r�b�:�>b���z#��}�Av��Wl&+A$�X&��K��Y�|HX�Ƌ/qex)N�>y>7 r�`����:��ED��%��W��X>�U��qm�TudP�}|�[zw��SB�t�5����._������"v�:b���ĝ�k�d��%b�~ϛr�����Ey���2�i,(~�nA�V�C���0GT���EF����H9��������fߠ��P2|��2��fNC��,�;�.�7��BK'OQ�̙%��ʽ+n��	�WY��b�h�nC�&F5���3X���)~:�ɺ>M�#��Լ�ڌ��kL���5���'��[�,t/D��0�W��6A@u�s������Y��[䈄JX#����5Wrw�U-z\���*9p�O�ɒH�ʽ`e�{��[�Dh�������Wx�Cګ��; �3���; ��N���j��c������^���s�H�^7���%��ˎ|��h{t"��[~��t��KI>�[x����K#�i��x�����=�cX������y�e���@Y.��Jzz�ғ12��6� �z��	�me=}�0��\Jbm���A"�)��8Z���4�u$;���o�Y��ދZ�h��?�/)e`��T�U�ޑ;�A�HҌ�a�����Du��6<��L�CF�������H�/���仡[�D�:�$��>�2��o����H^�~��T�><�7׶dF�1��(��ۉ"Rsp4��1�E6a*�.�##�P�JRݍU���^@�Q�$Na�f�8
��s�j��E �ߋx�{\�X&)��Ypy7�[�i#�ƴ%��[�� ?5F�W�}V��}&t��GŬ�|üSU���얾��?y��5R��ēg�۽����YW}"�����[�Ve:�:ىg�h���>�)��P\��K�	�=�l������3��S�c�z{Hț:���I	�X+ 8��ǆ{�ǖq?E㟄ϟI�D�7���adԨ��d���,U�����l�|i��+�G�'�nv��4�5����RZ���;wR�aXBĊ՘����G�c��h��"�P
����eXI�/����.u�m��cFm=�r�!��Ǥ�,���$/KK�UZ��f㐒z���=�8t}m� ?ȫ�PPk}-��+W��j��5�}.�ڤ��D`א�ʷˈ"���@��2�oԤ��qwQ����T�ҧ4D�Z�or0ҡo�k(�c$R�vc�OKZ�X�w@p1����`�h�@��
D`[�x��������Fg�f�f7v}Ym�	���/'�Jd��?X~w��v�P����<lu�m)���Y.�qlȚޅ��O�����
�{U�#����5`gI��Q�&R�`�³嫾��߃�����2C뚊2��'s�����޻1ڲ�'�c���M��/+�U%&c`�ZzNڽ�g(3�oN[/�X��e���Mq:��M���Q��&��}R���o�Po=�� I^�m�z�����LL�1"&^�YmÆe��m�65G�A���w���K��;\i���_,�c��M%�߾t �$b�0�{���WG�x��m��Xb����9�7�dR��~���8 ��EJ����*���m?��]!������Cs8�	�;�w��V��Ny��2/\�L�0�^�
����[xJ��1U�/��A �ߤ"$���2Z؛���+��{_�
dI|ß:��2Q7:!c0�7QϨX�:�:�LI1���ּ|ؼ�0=8�7Suw����f�T�fAU�Z���VyJF~3���C�;���>�'�6%4ܬ�^3���$�=�Z._�����M'�|M�]���	hOJ6��̫�� wG`��7"�l$�:鍏��O(������ ��/k`��e�V���?v�?Ή`�r���.F^���bD`�3�|�K��fB$�gn����_�x}>�~Zi�>iE���������Y�q���9=EFB�k3��w �}����lD��tW��ݟ�Sk����vKd�j�s����������C�L�� ���h���M��a$`��~}Қu����ֵ�2�%�����G2�(Z���dɿ����~*�1�e�W�	|h��Aׂ��M�?QW},[ڰ�T|g�t+�7��5_al�}"��5�3-�������#x�ƺ��e���)�Mu���c������X������ſ_��褣��Y鯁L��Bm��@�:~�w@�j����04/��r�; ��3)��Ǵ]2ge-d���g:Lz�1rzf,I򱓳C�s�%��OI���-���v��P�6% Z�ک�����1�0�L��\��{7%�+{�����-��߬eM�Q�A*ر��.о.R�+�cPQ��R�#4ckO�N0`�FP���K��7Bn=�_Əa����Y�� U��2��3�y�w�/��}suOH��5�9pݛ�4w�����w�u$wDݴ;�?a�qh�9����J��K��������/��t+٪&��+�_�u\K�};���m�L,��r����b���~v���8HL��f�Q\ܬ&Ia��J������UiX��U��,�tὬ�۪�T���_��`/_9c�Y_�):#���w WcS��ȣ�w��:�atN�|(�m��̛ܸh��?��%k�I,��X�(��A�c[��^�I�a|�_��~^��l%۵ ��İ�A���N�w���7S)��w��l��h��E,�aZ�������T߻���}nF�`���&�P:BP�X*����DW~�~<���h�6y`��=��g�>˷�R��r��tب��QId5!�?����>��D#�S��Y��DsHK�~�pЖ�ɒ����\�͇���ۅu;��v� ���G��&��o�5�n���|�f��t�
��c~"1�>���x𔖧�6�⥿&C�,k�/:�h�ۑ~'٭���U�[�E��,�ؽ�R�J�1���~�G ��K��)��VK���e�J��.֏�ˏ��s�L,QA���_�[�]Z+���JC�{�t9�ݝ<V�?��fS~�s� �^-��y�7�ٵ��
R�n֙*��QZ�?j�,P�߭�o۠�;/�8�
��Ա~<����8r��&��ue��i¼d��	�O4n�g�?�/����ì4��)�*�.'S*Y����R�ʞ�\���B��C{�cB�w���C
�J(�c\2�����P��h��`��J�8 �k{^������r�$D9���	+�6�����.���t��g�A���!O��(0ĬM�ǚ�P�$�}���0HRb��x�tcIE�/Ӗ����;�d���V?Sz��<�
&�˶x�)�Xx[E ��Vط�m�������'���� e��L�W�$w(`1\\��'���y�N���cEM���nj�e����L�"Z鉉p����e�#R�V� �l
�Ƴ|`�m��X�'�S����H�ᨿ�P��G������q�~dk�\t�eaO+ᤕ��E�&��Z;�!�3�)M�K�Nt�������7�?Z�&X�	_����	�?;�}�`��P�i���UQ��c�E,�Y��L��ে����'�a��(1��)�Eb���Xu75u�W���#��w�ӽ�"Ƚ��yv�(u?�l3}�\.���P�͝�|��7O���x�����<������ �ou7��@����*W����G2��rr�A�*���f��s]_�}!�H��c��z��'Thd)�㐮7Z�Xc;B^��C)�4��'[�g�m�q�7K0�4�HW�_��j�'��jX�����q���{>���B��f��r��orF�neR"m�vT$�3�b'�a��6��;O[��IS;� ����[Ԅs*8�3��.�ץ������^�ǈ0?��!��X]�ڈ�lɳhf`�^AE��	��U�w�v��*���ݾ�S��>퉶��Xg`$lm9�H$}J�� ������We����b��<��Tho�Z�ĺ�v������M�볅��a	��X��+e�*���n�4���R������\Xi�"���~�؝����K�J�������yA��b^����jq(�y�KیP��;�[j�C�!*���p�b��P�1�
=pB(��q������pz#��VL�Nb�u�ؤ���`.�FIs���[��;���-63&���K��}�c�c@R��r�����N��N�U���yE���9m����H�c�s⾀��݃q���)��;���@9�;�=���@�������(���cl�L(�ndd�S��7+x?�峓-t�������oQ����Ԧ3�b�g�ֈ��
�dh�n�]-SQ�wAb®ۇP{�W��y�m/3�sڧ�i��M�叄�_�d�j��8����&�	T���'�Z�^������<w6��p��͂#9-�^Q�-�E��"0���b���%�[�z2�w @=��q����3,1\	Ԕ����r����f�R@O|��?Z�gC�5�?=�W����B�%������jO#-#ź��K���f��Jse[ch
��P���mlg��M$U�!{e�#�(���k1�]�;�k�����rAºS�f"]2���QE Ȟ8ei�_��O��ָ�_�DV/9��s�n0��� 2��tsӣ��.��D71A���j&�1��iR��]����w�靜����'524�=�"�j��	GsO�ٔ��[�=�k���T��A���ŜY7������Ʀ�����!7�f4xB���~���P��t�Lz��?�m ��S��m��R�4�Xf�u���[bFJ@u8����fu��e�|���޼Klj��X����n�%�-�2M�z�}e���Tsv{HV9�$�x�B�����o�3
�2�73�*�ОK�1=�_�+# ��d��2"�%������Z��F�I����ھ&vU�jh���'Ž���3�= {���S�'��:�S/��(�̞�1g����>�#�fC�}��X��_�� �%�������Ծ��3��S��]�'r�/&�5Ŀ+h/���+{j��V����5b|���lnC�^wb+!�6�@�z�4���Z'��lD:;���h�Ԭ��fP)>,�}蒵\kZ�|���PG7��t�!��A����ݖ'�bu�}�>���h�I�9���`QE��sdYR2�K
M���?��Z�N�����4��;�S��#\1�s�	�����O�ⶻ�5o��w$��9<���d�h���J��/x�a,�f��3���R�?��nK�k���)Ȅ��ǻ�;:'���}m��8�<��NHP�����N�J#�����E�ϕΌ�@�2�j��Vش���jԶگ-_�0F�i�hپ�3����x�;�.�� =yj{�v�y�kM������>K�|�˿x��i8��y�<"3�:�V�jx4j.�x���M���c�k����`	6��G��~�5�S��j�2�XÆ,��v���ccsi�f��7k��Yo�6����Wk����[���a(��.vi�g�|ƚ�qyHg���'��l�;�W�;��|S#Q�Y0k���s}Nʵ!U)0��{����_��t$��	>�- �Q���u
�mM�վiX���5J�'ښ����8�n.R6��ds����ZqH�k�veM�%Ax�s�?Ċ�A��Xc}���F�-��E���)˥�/F�Z���C�ʴ}�DC|�čP�b����l,�@5e��'ߪ��<��-e5�����\��д:����o�;S���!<��^d�����F�r*����[�Hsk*��?�L͔��M�ɂ<���[{����ruc�I�rL}�5r":d"�޽d��t5�2�,R�ԍ�y���<��4�9��{5;غ�	�Ŀnk��}�νJ��|ؤ���)I��O�`�[3�vk�17;B`R��2u�k���i�&[�ܠ?Q{��G8y����$��6ɶ�"��A���ӟ���"��W��dc����R:xi�B��w /��K��Ӏ��q��r��,%����t�m���С�ڴCf�ɸ�
�w�P�rn�`fQ[�e�*
�kxf�7;逷b��	1y����|Ro��2`�mް��^?��}�?|���K �ަ
��-�����H���Ţ�W� ,��u��V*�ۀ��Ԣެgш:��9��>v��;����E��!26J����� ��������t�~�`���6\E�h*j�~��c��lKU���}8y��Z��\F��� �����&�K��yGµh��F(>ߒ���u�#�ޡ���Ҧ�៍1�_UYi)/�Dm����w2�&I�w�y���y�0��n�έ� ��+�릇T[L�N)�����{�~���W~bA-�'��W�'�Ƹ�Ѥ���K�9��<��$��XWf�E���}"?�6lYom�� &|P�S�-_����F�%��r�ǜdc��E�W��&����tRm]�s)=>g��ry��1���V`��<r���w��s���9_U���t��H,��72'@fox߸=A���l�c�4�Q�9c��ڦV��X��<��W�ޤZq0wʡ�Y��l�E!57�Ny޷h<Q��b��Z�����z�|�{��������w����\a�o��)8����$��:)�n�t��i著�#ʳ?';�&���x_��J`�[^���
�s���~'�
Ë�-G�m.U�Y��Il�\������ls��0��L����ҐT���d�F�\���-j�f`���r�]IM��k�[��L�?�k�J(��S	;���d-2`~:�������9L�?�L�?9o$a�����)l�ITL�IW��o*����%a�מ�1qa�; I]�O;l���3���w@�kú~Í�cw��I���
s[��Z�L4$F��Qi^+��/�Od��n���ե�-/��{����zT����[x:���+S8�E��� nP�B���b?�t|��F��a��{�����K)��v��:B"�}\�K�`�AcR��z�+���/�+
5�#�/�$�p��W��n��+�O�_m�	v'��;�I��`ĉ.N%�q���]�|�8tku,<�6ˏm\	�ɝ��g���ڲD�sZ�WR(F�K���#��'㕁I�#��K޺u����N)t��W����5��Ų��b�&���!a:�t��_W7��b��%k(��ߔ��l�7ٷ>�C�Q�u�����kJ���Sˮ����N�b_A+w�+� Q�,��&�W�=f�,��1����f�����$�G	㺦1_�B�D�D9}�9M[�'��5��~��������0=�n����=�\��o����K�����g}�S�������߇
�L|z�<Z8]�~k����.�Ƈ���5WD6Q�Obm}���4C]�܈�N-.w_G�q����Ϙ@`N�1�x�4}j�a�B ��^�[q�/�7��V�'��+w/&���Xcӛ?p0�b$��[/O\���M~�p'lU�; 2o�b�޿��D2�����Œ��kng~Х k��ڇQj��4wԖ�Z3�"ݧ|p�)� Ų�0���s�4� �kY*��#M����*����?���^p�l킥a�%(�Vx_{g���.G��G�1�_�:���h�O�NB]G�X�i���/�P�[���1�1��ל��&h���JcS�E�䇙�.�u=l۲e�Z� ������a���
�v�� ����ӹ@p�*o�:7T!/���@�{���oqm�]4@edE�.��^��d�˜6]C����i��#����.44��f�ɳ�Ҫ�8s���8�����w4˅7x�\�_P�u��F�8��Z��KI�"����_���\�v���낏�.�d?Ij��W��sҵ���ܞ���y[{���#�x"���e�\W��W�f%wZ{�&��K�+� 0�hG�xs�$f��uWr��Z*���+�@�ńI@�+"y=�DS
���,��ޡ?�&E�I�������q ��7/�X\F�65�|њI�Dy�_�1(eh� e�ɤS���}H��2G��&����wwH7�dOɾ���ק蓏�_*:Dc)x�w�_?�]�t����؉ꏉҋ\��ՃWB5�+̺gQHv����wor�?Y��^�A��\�'�\Y�r	�E����l��o	�ds�R��)��>&�.��-У:��C��PvT����Ո�./�״�闘Gn�7�k��>�����y�ѻ�w�u?%}A����Y�-�,�1�y��L���)bfT��:�9^�[7�4�/en,�W�l!6H�wk�ߓ~��Y� �x�>e��)Q��Ӥd' �|Ʋk�<T!ߒ c�������UZ���ԚKm��>��k|���*Z���i
^^���0N|�-r��[_�B�K �qC�yA�[���C����

;�l��VMY�z/�/z������p�	��qy��
$�����pf��e�XQD��˹_D������$�����La[���J�z��>~���60j8�h�SWo#��2���ȇ�-�{����;�ڭ�y��Ӵ��r��\v0H�λ^CC���`��5Z��˔���HC��G��跦�ۤ�e�@�B�ͨ�Œq���*�3f+s�(>��(\if�E�摡�5s�zaVh���F]	���mj������\��X�f>vM��<�x���"���#Qل����áDa��˹������w��3uK�!b^ŁN$�W����KQ4�����p}����t�l�� ���
 ���\tgke[���wI��ïx*�MB:[#�|eO^Ϧ�|�9�(j^f��cmkg�o�ؐ�_�xQ�����L7YDwA�4n	��Yi2y�������φ�	d���nK,���y��n��U]/�iP`J�Q/��/xD
Of3I�>�XM8�զ3M�D���?�t޴n�2�w<����y����e�1������Q��s�C�a2��NFwl\׷IՔ�>|�^��V��^�8��@)*{�]P	\m}��}�_a���.D�}'#�H��ӸݑF��f*�a��)��6͎����0��_�y!5�3\������X�����*�w~ͱ5��~�qjd���h]����l̦��m�'E?{��+0�7/��->�o�D�(\G�G!���r��� �F�YX�΃$%yֲ8��Վe;V�ؑ��3�Vr�}G�&	�O9���n@��]��*�3���� ��W!�b����a���{_�_��P4p=��r'��e��f�Ծ!w��^)���p}���n�-䄊!q3տ��CvӜu?Q�S9�7S��f�����g�L�쪀��"x^Ws�r��m ����sK�nŹ�O���;�6�>����_m,�}�d���������Qq����.����\��IQ�yq�*�2'HY]��S��Q/?N��DR��
��2Ȃ��l����k�2��any���Z�Y�9G�Ǫ�+�*�z�}2ץ���fr��x�����Ͽ-��'��/�O�*Um��	�ՊRAM����n�{�i���%�%���b��z���i��RM�� a�X����y���{6<ً%.ZOu�cu��u�>0R�N���٨�#ǸƔ��Olq� P9����Z(���X}x-F	M$�U��N%F�%��褭��Ǔ���#��3Qm�V�ގ��3a�1��b�r��f�j���U_�u ~�zC�Lsи����
�P�R���r]�>�h�։��1F�'�(n&�zs��+UG���6���~!Y]^�6�ۤn��+m����=�*�O��r�,�	tds�,��cD�ԙ��";�5���^l���V�Г�Qj�{�(���\����LUu++ �����2-!9���T-8,d_w�Yb�SV�Uo��0�S�f��X��A��[M ��w��;��������km��g̊����!Q�]C�t��{c���Vú3Q#J�%CO��b3��y3� o~`���Aҹ�[A���u~�5�VV7~�K9K1��BU� lA���2���}��q��g��+�.��sTU%����Ԝ��h�ꝁ���NK~h��+���݈��[����%�tI�3��Ɋ,��!p�h�ڙ|a���u-H▚���@2v���0�+�'� Mn�R����5�ܸ|�v��F�c
^��I����U��i�h�+U�HP�Nz|�-�:̜��[�[�� 4��@��O��� {��/ː���2��ֶ�2���F#�p�?M����O�:�j>6�f�e�}MϾ��{�8GX5rF ��^;���#��D�e�X���E9B<�k�U���!�Ҝ���ʔ�l"#�	%�v�������X�=xX�_�X�
[\�Gh��#�y�ʫ�8�UR��E$�'Wq�e���umŵ�s����=�>|	hMXK�&ͷ����)�/:����.H�9���a��V6�Gl&�1Ө�>3��U��h�5^$��9��k���z7^F�	����֟�{͹>u8�ʿ�K����z�P��)�C?��Nwُ���������*ꋒA�qM��>�/��^�Oe�뽩>V�b��Cg��2� �<��6�����5B���kA�M�=�LR�f�_Lx�t�fDO�\V�:�llc(o�$�|���7�,2�x)���S9l�:��Wn�.l�qV��JjA�|�k�x��֖�X���|�1wwb��\��,���	zw	̠>&D��
��tOd����N�� մل�E�/@���L��x#3��]l�@AQL&�mu�F�X�{��P\��ԭ+���ZE��W���ƍK�a�MU,��qDC���z��y�w��{��|���f��GUQx�OOI%�$}���;��߾�!N7��Hj>l�T'������ã���J
�N��Tz/��FR7�]�&]���n�h����*�]�0�q]K�l6xiΙo*��b�-;y״�8�X��e�d������?K���vX^�n"�u�0F��7�������.g��Qe�����|^���/4�yۘ9�����EC��j������0��9����4�U�;���p~~ݯc�'����ׯ}+'�9�;�g7OZY�y𳻽_Rohjq�JF���B�E�!ͻ���۱�*���|�ߢ`����A�5�I�����F\e��o���z7�������V���]{�}B
<�����`�L��j�Y����_Aw�2���a�_�z���J�wM&-�[��ix��{�w{xX)�6uK���s@�,���b��v)�H�N�������uF������騢��u�h�UJb��I�ɕ�S�X��(g˾�'r�B8�B��ll,���ᐡ{����3>��/W˙��y���l�O�9�����%���r�Hj�O�'��m�3�gyt�o�du��.���H9]����ԀD�Ko�B6��~?fk��1K���YM��;`x$!��CW�)Z^O���^� @Ūe	������Kj!/ŗw�����`�r�&�L��s7G`8Ny�	̳��ş%�B�������nA_Z�5zVh:�+�������K�j��h�]"L�k*�?�%<�ݳ�TO�۷U]��c�AP�[WwG6�R�6��J������$#c�F�S%����F�����z��֘Uj��^���.7>�1Rv�[���/\�vzًD�%Z��bI�*۔f(�%�xZ�KB�T�*~�!��bp��F-��ޑy˺4�0���֞�?�t<��*��|4o����!�5)����7�/�(�iI�Bu��>ւ�ϚC�5���޴u���Y]�����D�m�B;|1��K�i�/��n��`	���\���C[��sw\C��k �����%�YP���
�8�a��Զ�Rmz��)���
�V�K_�A��9����B��a']�F9��L�����h��L��j�s"�L��h��m����v�YX0䬂
j����¨b4�����J=4�&�O�Q�vC�C�4N Q�^�䝮R$����-/�/\fvh��7<����S@ܫySf@¢���7k�B�x�$��L]��J4^�T(x��H��q8������c��銼����32Sxxٹr��t�9��p(/'j���7t��ҍu���(�jӒk9��&QA�ʉ��F{:�$T�i�/$?Y�f:�m���G���o/LUu�#n�f�N)=r��q&{o�*ՠ��ii �>^���:�,��,�H:(a���t�����B�hO�SKo�di���Yi���W2T9#���:����0��2��?3/]�i?�;&XR�dű0�(��qU�<��onM��(�R�c]����ͳ���wƩ�HE��;���[�y4�MS��)xd@C�r9�} ������������a4��bʸL�;�f�(ʱ�$�D9H:����Ef���Y�ZB�,V�u���mq��a��׉ݭ�O�2u'��eq�e2�Q���=Δ��B0�|O����¤nV)��f��գ��$�/��M;��Ƒr����e�Eo_Δ�γ6������!?L� ��կN�_$�31��Z1�u�] �d �_�7�v��b ۀ1z�+#C�6=C�eyk;"6g��
U��'�Ӟ�ڬ���a�3��� ��N@�$�r+�]:��1F��EӑY�x{���ԃTW��VK�5E_[	��]����\�s�8Z_"`G��HԲ����IP�!�@��~����&��s�0J�C����:��1f�_*��H@����UU5����ƕ�Uhh'�l�Fg�1(BtcB>�Ɇ��������q�@&+[���0�oN��_��Lm\ۤ�ϺyN4b��[��q�"��IX��:YQO�8�G��@�'�d���������ϙ�
��O�F:m9�\+�z�{��>�Ǡ���3��{fu7gI����-��U�ݵbSé��-��}����4ud�*ezA�O���G�[�E���K�� �)ݍ�ұt�t| I��\:�c���P�AjIA:�c��������ݹ5s��q����̹��l�$gœ�[$��-�K땖"5�D���7=p��e�����������ZvA���ٷ���k:_]3�<#ܬWƫ��rq6�c'�r��ҿ)���`��[��BSr�Ti��c ��-I���:���� ��%��>����v�Cn����A�d�4[��[1gX��H�%�9r|��E��ce�yN��5Jz�~1*Nx���Gi�V��o��~P�(ʉ��<<D�Q��V`�7T��Lt�7}z��R�Ǎh4��'��c���A���c{R�@�KQ�	�8u�L�51'�7�����<�%,�mA~�j.�{/Y2��1x�8��d�]*{�ʢ
��f�v�Fx���®�Q��t�xe�V	 E�m:~�ʉ0���[�q�G��$�)����{�n��"	,�촵/2޴n���,%:_����l�"?[��a;p���/`��h��¾�~Aϸ��֩�?V���Ę2WPmy�6��T$G��]ꪉ)M�H�{������el ��n+*n>�ѓ�	���m6�qv��\�pu'0��f�D�׮����d���Q�G�윃���A���UFUF�lRa=��J�2����ř��u�O��
�?Rp��N�+�U�wf�jeh�r�7��[����d\�,��(Kv���l��F�L��6"�~��';�P��ga_CU�*��2yy�r|�t�c4&Lݺ}�An�`&����;���'!k��F	2�`�o�Z�P��	���eV�V�1��:o�o7�E69�~��喤��ݴ�h�tO�}�g�0���5�b��8��Jڻ��ZI��q@��-Ͻ��Ϋpl�]#�/�D�������R�'7�����x��h��F�����\4��g�n��Gg��(6�F��H����:�E�/�W��R>���QٕGtsI��-|���9o����4yc˳�o�$J?m�1�� k�I��W��]����4_�v���I�P�F�����>��"��9��~�>��縉��c��Y����{�~hG<���Ӫ�p;xI���7���֊e��3D��+wXب��4�t�CMi���FU��;�j�g3��s�7ѭc�K��^x"���;1��H,��R�&�oo�\x��Lӳމ*�l�T=L��EC��힒>�L/m�W���ɾ
���Ǻ��u�u�[GQAg
�U��"yd��M��X��G(��ɶf��b(�V٩�����t ��/o���r���ߦ�6��{������e��2^�u�h�a����KR� ��rA�F�.�d����Ɖ n��A��ydÕ/�a>?f�{��&V|U����z��/��x�e�}�͋��/Lx<����p���Э���*�:\�(����/�\�E�N9���x~y�VO��aq�C�a�s^w�;2�^_ R06�u_�/8��������~Bk�d��J�����h��<þ�/���4B�h�\�⵵$]�<�m���+@��؉���r��7�J=NM�$�tE{S��������!E�Yg�$j�⣧�y�&H�e��v��|� ���_��P�*�"��A`H��� 3�G��G��	Ml\����z�*�C��q�a��i���^���X�[�N�B����6�B�:�j�=���t����9����Em�Q�	��-�2���#����;�I�%uPOOk�b�aAhY� ^%�&|L���������o�4�9`�Ta�Rί� ��fLd�
0Q��O)�9��K]�
���@D�=}zl�F�8<�1X���_RUr&2���r_3R�U%J�J�����ʦ�	5�ן��y=��J8:�K����{^o-�t�/�\Y�h�7�W�8��� �x;|��8�<�\k�R[��R�S6�C̜��!'�����8��b_ F�5��QS;¿�(��i�h�ѓ�C��?���	n_���x)�����/ʿ�0�-6����>�-�5I��o|v���t�7d�H1JП�p��'��'b(e��_O8��g-�[J���_����=�W�� RG�W��1�N+�����2ޛ�x����VGr�/]��S!k�3汦�C�l�/^"B�SS�vZf5=�+|S���p>�����)]�3�$9��S�D?u��Z��D&�F��C�z���l�Zg�6�熗��c8ܢ��#/Qz^ �[g�b��]m|:��X� ܙ�1Ԗ����6���>~�
v��?�:�(��1�;����>�w��4d�-A�鶯��)y" *�����?l����b�9�����-x��߫G�|d�Bd�~��,���#s*���V^�����l�}�q�p����*o�cׅ�[��:������[ͫņ��x��4�ҍ�<Є��[�2�W=�0���/��Z:a���F6�M��<����.��P}�r�_*��设N���+���үY��:_5B�xͼ�Fu���V�u]?��*j�<ͼ��#8�C��婐�zX���ء���o� =h�'�2> �"�nM�b�]����t|*�x�Ĉ��1�����!��;��%Z	�V7��6�6�~:��ux(�{�}�z��<�i#�6�FW��9��m��P:�\ ~&�[( eT��Ԫ��V�f� ��;�gw+�K?�� D���	kgN�Rd����w8i�z�RZ ��C�<�����L�:Uj�NG��Qa�Pl,��J야\�m��А���~~}x(�sO�T�����L@-*���nk])��۟`��@A� |#�d3���`���V�TB<f%I�Կ��ַ�-.l�#��_$�]]vIyEq,�ؔ������>���=d��!��*�f}�zY�����=
	���3�B�� �-�קGnl�s_MZ��̉x���^�:}�%�NK�/� F�↾֥�m,u#m6�m:�T T9� T,"$�e��c�W�U�M��)IIQ\Vy$�>*�a+j/��ϼ
KA��h"�����0%�t�eba*Y2�[f
*J竭]�}}X!@q�_,o�2������{5`��.��a\���AR���Z����m��=��о~}��ۧlG��E�o�'�(;����jB�U��.�~!�O�F�� As~Pa�0v��m��Z�0��B �r�.�deQhh��U ۿ�l����ҙ�P�ʟ�.��v���4?����fn���M�N���\���bG�L��EwU��'*)~TYԖ��=)w!�SbŹ!�91���u�i��e�AZ���#ݸ���fۏ�s�%H���$��F���3i{�[��36\����(����4n�Z��f�q�$��!@>n˾#Ⱊ��������%��-�%��ji�WK���36��jt��R�,���܋R	A�^���/�o����7�g��x�ښ�YX����#�Pz�%��C�L��R�T��LL��.X���뫈��,~׺���d@�^��*���#�ڔ�MhP�[ /�J@^��C�WB�W%&p�������8F&�*����۝��+]g։C�KK_��nPQW�cC�?�Ƃ2�LY�j�;��w����GDl������,ce��x~Vk�T��+��3_�6���|���)�����w�c���dhD%gp`#�j����\�/�g�Mi��J�HB��N�]�?2�����?���� e�p� �w�u{����"��ϲE�I�11�K��u�1���ҹ3}�m犾.�f��:�n��hb��C:��n��nт�=w�s�qh�35Ƈʝ��m��,�qD�� L��}iHґ����3��Z)鼵0M�O�����$wz�#-����xi�\��3,zJG�*�Bd_e�d~(���<' ��zB�k?+�g]Hp,՞+T�.�R��f;��8�h�a���b�xP��`J�c�y�}M�<Ovj�8-/�F���8���.����NmUe�-%.se��K���얞���.~4`��`���IS�Fdg�>uЭY��kkx�JM�ӷ�z�e^�nGhjR����l�B�K�UiY�RW-wk��&���!�K���^���E�{����]��*�B�P�"�}�	jq��� �ʗ۷7D1����}!�z�,%\��`A8's��Ӫؽ5�u`��5��Fѡ�	��F�N�s.���x[��C�r#�(�ۤ��?*�ݏ��W�_���5��V���f�՗��� v|`Nգ��ki�����7%�����x+\�p)�����G~FVK3�.jmyN��^�wR2N�����B��;u�� ^�܃M��c�7�M>YiQu�A���Q�������ju)�N����>]�� +<��ہ�h�~���� f~���ܩ�q�P*ޜ�J�%��%$������v���"���U�Y���r�Z����{�r�9�k����l�����%��ž"l����%���$�=���ɉdgB��\9f��2��T�S��:�l��#p����NI�5J�Z�@|"���nז�9�bd�����8}g����Q����!U�TE@���Tƥ��B�o��N���� �7K�ͤ�8�3�K��2d��(��P��фB5��D�7���B��8p1ľ� �"�E�/ ���r4�
REK�A�O ���@���-9Li�Ś���]�ժ�8���@�����ӱ��M�Y���0</���ؕ�C��#�X�שȿG�D9�_������;A�O��uĐ��_ҩ�K�1E��iS�؅���x5���>.��0��M�_�9�c�@ǖ۸�ė!�zXu����W�(7OA���ڝ#S}�Zp�g�o�E�:=3��s��X�g���5�u%��&�3p�8���G���x�j����r5;5
�����~�����"�l�Pa�a��('M��`�"�J��`,V��@+�$�d��iѴ�^�_�[���"�i��̉69k��=Oyn����%L�)x�<X-��n���I�ET�/^�j&�>�d)!"�jB�a)���`����B�,���T���ؕ��}�����ɑ�F�l/�Dh��]�iH!%�Mޓ�sB?� e9ފ		R��؂�oW.)�a�r�y����/t'X�U�?1���t�(В]��`�>Q��ĕ�d"ﯞk��*q�	���I�h�q>c��K.!rr��g�3�4t�K�mA��7��!��LvB��Zz�Q���ԳF��h���(�{��}�r+l�z�-5����	/ *�/�/ ��͆���q,�vobDf�@�8�O#�\���-~r��f�D��t�4-�^}m�}|�����|B�V^*�&�x���!�-�ɠ�v�rN�Ƃ�rG�4�.E&Z0���P������j�������ٷ
8N%,!P��� T1[;V�A�����2F�Ω*~5������حL�!�UI��"���|����1/9�����zO7�.�U��$���
j���BSh �O�ǻ����Ef��ᜧix���\y�u����j6�����hEDĝٲ��=�ע�t{�U6%6��\�v��-�s6-�?�.�r��x]�V�ɣEB?���\��+V�Z���L���r�Ԫ�Lf&��N.i�D=�?��tGq�}|֔�o��q�pŰ����1�&��,]���e|t2R��!��~+"݅ťd��*��)B�8P�������=�����JQPSu���������ϓ��4�SJ=)��X���G���eť�:z6�_yH�%��r�5�#]�R�aُ�dRHiȩ��j]�b~�@7q0"���̣�qM�C#�W���B��ZG9-0b�{�o�g��L��<�c�n�_S�2���JO,<�X=i���T��^�6L��B�a�Z[�������S��$OHb�tkƵS�շ���E?��'��i�WXz:�;GX��'�,�H�����h��	 �&d$�۳�g�vpV�x�Qt�n����v���*C��t�\�3�۟U9����ǒ=��+�`�-��)�,�,�����p>�����m�6Ƽ�D�}�S�S�T`#ۡh��C�"#��H#���m$yV�8���:1MO��|�Bvo�9�8W�d�$����벥DJ��z�VǞ�B��g94�-r��X�G#gH�x �6FV��st�;
�"ü80f:�12�PltY�.�XT�0b˩
<�W߮����S,0r�Oǖ���7a"����l�#V��4���������vS%��c�E�m���o� ӽ=�;>[o�o����O�ʺV�������츭��/t_�~JIp�+���#ezs�e��W#tQ\�6��\��G�(9��0�Q�`���.�.�⠢�+k�)�%�c�p��pq�һ��]�op%|S�m�靧�K�[]��S9���Jg�#��U~>�]Gh ���s�����S��r�]���"|d��|f�
@��{E���)CK[M�"KV��pqȣ�E���a �`a(��j/n��߶�U�L!��!�%�a�ۢ[�����g�o:$�g�o���8\y �A�.[��*��L���������>�FVR��p�8�9x��+Kv���a)PA�lld�$��8�ۓ)W�p���g[��q�����-#�꺌�)G�������y��7�8�/�6�؊-V��ָ�7���)�t���6k� įn(�g�B�9p�j���q�ޖy��%�WQ�F�O>A��E�y1rE����nh�V����\�$c��.?a���@*O�^cy�u�Լ��Q?��J���c�����oCt܀ ��U{��є��(�T�e��>�~�S�J��D�½N�'�0�e��-cۥ������<֊�$z�V���X#._1�_�\Un�d{ة�U���ݙ�Wy>ը�����HQ��A��� ����,��W/��v��ƫ�����O�,Ǹ��|%�Q_ f�t�ޡk�I�� �k' ����c��id���ЩX����0cQNqz~/���k�&Pi�l�WG_�d�u|����A4xv[9{�\�A�;!���(*$���C��[��7dJ[|�if�|�kE.핝�If<[�����;߽�<yxѓ���� XM�]���|���������<ϛ#S?�)YGCg���V呣�,�)��e��#��Eym���ՉT�������1�uV݈ސ����[_
?�����:��pN��u�-� �|�Nk&�����N6|.���� �ng���r9I�Ky���kه�+Z��F�Ϯ��e���I˿Xb�uF��1�e͂V��~�mwiI��Z����>L�+��~�Glz)��i���yZ!�= �^L�[�D���������x���k�z'���B����j�v�2�cup���y��+�z��
�8+_;A9�kP�8���0	�7��9�qr�4q�dt�Ϡ��Ӂ�"��8��¯��b�6'�V?ǁ����;�0�N��-�3Ua0���hN��#���-:�r��+���8(�n���`�C��Y���6��\l޼���(�!<<K���$�6�(h��j��.B8�]�[U�7�跄���2!~�w.ʔ�wh�6�8rJ9��&h�l��)��A��N�Drb	��ހN�7_c�HR�|PҖ�����i}���Jk�R@���[ͻ�q/��Nq�7i�@c���<���U>�G��ZqEI!�>U.]w���deJ�ɐ�A���#(��4�4��8{�A�W=��~�_��柌+�������(�:��T�N�Y����W��>��E�u1�\F=:H�]�{!Mw?�����z�*4�d��MA{��5ִ-t޿<�;��idf�W�=m�-��?��8/T����zf��Э5/�׉j��:�W=��0�������6-�p�5Z��o�g�:�0�)�>�#C��Z���s�/Mq��_�n��~վ^^�/Z}���BΘ��Cq�N�����M0�W�W�ߌ�k ���KZ�#��k���<u`^-_7;:I�p�(�3���4��ĵ �B!����t�E$�`���Z�[(~�̏o��2�@��ʛk9�q_���G^�L�_�wxY���ج���9l��z&�%g,����_X�8V8f�E�9~��H��t��ݓJR6�<X=�-�����&g�^E��5�@��v$�����Ƭ-�.7I��Gv2���.P���Q�w�;�8߾���3��mg��j<{_�����γ�4��Ƶ��49�z6^k�
����ʳ�Sj��ҜnW\o��ݐ�)�HE�bXs�}����GZ�+-�ʈ�oԶ��~5�`�M~�cs�Ϋc�/�j�$��p���H`�;�x;,�_[z���^�d�ە��c`��Yg~����5��!0�@⳩��t%>�X���T�pA�}�Ç?-��v�@�/n���P{$8�Yr�<XH['¥%|y�|����X��"�SjΡ��W�wɪ�4��G����=5ƃUO^ ��ڢ�p|`�~�Q*ę�$�iN���նēq��HzE.A�W\4B]��fª���S�����r#�ґ��Y~j!�(}6ڮF���Ǐ�|����G�W��5��Z<�}F�*��@RkA����]\\;@��ph�����6p��T��+-?�av>J�t��s!w/� ܗ����4)"��ji��Գ����vϙdƘ�}[�x�ӟ�� 3p��9Sy��E����_���ӆ�u�+g��#鵿�\*����|��S��IH۔Z�)F{3/*�oWS\�/r��@2���pc����1{��>�ڠ�z�����{��o�춯� �Yy����ⵌư7AO3��^���n|�)��?���v���.���>m��}0�PCw`y�h��ׁC�ŷY;�CJ���ңl�$�@cR�Fb�����R��з��*��,�d�|����x䀜#�5�Fqe�iYB���xx+�YJ]WgɈ�r���.���:~� ��)�����!Ԑ�#p1�sH���2��z�Q!��P)5���GTfr�;�&����0��~r��������U}Ӣ��X1�������pud�zA��n	hqye���/�7��x������kA,�yا�<&,�ڂ\WP�Gz��F����(���sj�|q�B�����O:^&��*���֜��D̾>rJ��0(z�j�:Ǻ��q�^�S���@m~�"��U~�v^E�SS07c˰��m�Te�_;"��+�X��#[�T �o�;��ϩQ޿�6���B��=ʾ�YuhX[Ӟ�'�^Χ�����u�h�X�m֌%�	�8�).RBS��Z�&ǑQs�6&y�G�ME�)y����e'�̱�T�2EB�Ǘ4�Nu��L$:z��|��n�<2�0�K�B�j�p#�Z��Bn׆� @����	�dv��k�fgT'�L��=��L���R���`�#11j�_�l�*e����8�����	�!�T��!��/R�=E�pM�6I�])Zlxwv۾��l�-���W$`�g|[�P��?���y0�L�{l�F��P�Ыo.��E����������',Y�� ��o^�s=�zMA��5�`J��~��Q9�Q*����4��@U��I�)�;�/����i�Eds$矋Ⱦ<|��KS��+d9L#�%��5�C/�r��E	;R~M
�0��e�8������"�ljov䠕J��������`T���d�����Ư~4fu��*���$�w�s���g	AhĦ����J�ߌ�<wbNF.��(9g�S;�DSU�v�M����rt'KYGXGUl�e5�=��Z)N���4���Y#���Q̰!:1~,=Rrm�߇��YS�K��P�c]���*}"$QaG���������9W��Vj����?U��\����������2���� �+����Ŋff�d��%�D��z��gd{}��*���B�����%�JL�Z�T��+Bǟ�[������!��O!�̲�Z-@�'ć�'�c��@�{-�_�|,k��m�5De8�0}ȇ@	F�1N8��aw�$r<B�u� �������,�~��/�W]�ɴ�W��@�m��1�Ͻn�h��	q����"���8��J�0���6uG��ĀNQ�Srxx���8Y���]d���T�c���X^L6��m91�}̊8��f>6�����W�4�mX/�6
`�S��Gz�]mxh��V��p<���=�*�obzI�{��"LW�������K-\����#� 1:ix@T7`���������&�gU�z����s�� �⊏����ƫ�45���ȫ�~�1Ű8�\]�Q�R*uHR����+�ؑZ���>J��f�Y�iDgYl��;Н�P�&>��3���� ��jS�½x]��c��b�����}]�fƂN�|����]g|�'N�ʬ:�Ö�,}�����(6ʃ���?978'!��LMA�ܾ�qr��f��d>	a�*?L�K���K�u�~�K^���e�7�6�<�Y�H�����*`�*�`��W��!�����T5hᦝR�b-�y;����F����$�	
Hׁ9��~���R}℃�{�xk�Jiv���S��!��
��4D�F�y�58�i��Ö�kk
X�o��{0�@�%��W�B�Z��[��x(�6�ϊ��n��bI�n�,ˤ�����m-� �A�c�n�����S��d�1����>�t\�&d��VF	����s=��e�.������a���ib���B䔪|���q�h��?�T�mA�^�sK���I�J+gWSz�H�>���N�:D I�0��PJL��H�~���ޅ��$��v����>�p����*ճ�ԇ�r���~�j��T�_=׍�]i�TQ��\$�z�
�Y@�g-C���Տ�Mr5�8#�o��"�Y���d���Yhi�`���2��,H�P�Z�:̳Fez/����/�Jy��=��4ª�}�f�.�Y}��|g�ܬ�Ml���bn nS��)E���}���@��ϔ������dǚ���D�I�����0lr�Tgw�J��E,6�ɛ��,"���_�8y���7�R�Չ��3���b�ՙW��4������F�-�ϺȰ�7�@�����5^��\�OS1Hs@d�5�Z'�VY�6�ݶ�PSQU8�Î�qM ܹ^�j�n�%j8����e.C�d5�m�g7Gak�x¡�*"��u��7etP��+��B�來�tV/e�~�l�S�\��dF�8���h�lsp4�T;95^��	��E�W��;���	Z]����}����I�
��OUT�]���p��;r�g'��gh0I()E1]���=��L��'u�Z^@��gh�LLe�U���w6��Ľv'��AbPI�*4��g*)j�ʿ-��QJ���
�������i
l�=���ِ�����1��*�QRz�}U`�~��� ����S�}�����"��o8MM��'��z��_#��oJ!�?|D`�P��j&5���7Z5�����58�����[�]E-�2��!�H5u�+��E�hE �8�3"����a�p+��f�Ot�o!�o�y�ַ^(i��6���l=�o��M;��sH�k�nW���=!�x�+���}�-H�S/�3s��&�ė[c�Aq1s�\��hi���*�A�0�%n�6S��{(ϭ[��N`���w��_)�Q3Y��Q�5�@L6�m�3�ʲ�CW*���@�:�(�.�;���܊��\o�݇n?�
��q����׾V���t�Q���Zz�:����������~���'x�w��_���e��]�P�i=b�+��%�΄^KX�����~���Д����t�_�|�{,��bX[���Ȕ�+5�S�9���//UN�VC����7�Cy�Ne�<&�P���f����k�,��jp���eA�6ײ}�pc iP�I�A馪�bǽ^e�'�z��<��Ad4c�O��ad߽q���Ԩ��^ �s�0{ %�H��<,���"7%mW��s[��x0�J�|��(��|{~��KGz(a�\=ۻ�+M՚ �~�u<EP�Z�.�-��,ߵ@�X���*�P ��O�'���uS:4~����
K�p;	k4xA�q`��ÝFEd�
=��۝c��͸Z%&��q�ʰ���|�m���U�e)t{�-Ha��U@�XF�}�0�Ɉ��g�3!%�F�r)���:�9�=����/]B�B&���hm,��L����
Ls�η�Xml�+t�`���u����D���������˦���u�eNU��W!PF�['Ǝɲ�y�W/ ���1����� >�����'i,��v/���
KeR�Itx�G�0AH�Ѩ�Z���@�s����[g�*ZS�
M���S��cxﯕo�RDK��Z �y���@u�^�j�O8i�N�-c�I���gM:E������q#9�О����=2O�� X��\�k�p��[�+�������++|���9m��g��zј�������=]��!띶��({��2����#�2�H�_������}	 �9%�t����[MS9�]Ky�<t���w�\H�}���ε�GP+�et��lP����W��V��,cӿ����V'0p!2Jk�P�	Ҙm�W�=fo���m�6J7v�~恝c��{��K��Hl�Z��g���ߕs.�G�QԊ$g��a����m[uvڛl�d��&�@?�n�5��v_��F�s��=`��7?�X ��%�Ɗ���L
iOZ�8B��Sσ@4�Z@����2����S�םc~��}�C���"_�װ�f����d�(��]Hs-d�W�.k��{/�*|YhI���"ۙ�'��5*OT�P�W���z����۟��Cf�����)�~Vb8׆.a#(�xW�;�ezB�����*ƈ����ʬ���$�&��F��d� ��%�����6�tSU)�7��E�)�(���8��#�.�4��W����E�k��}]�5�l����;5�����w�N�L@�yX�>��)
�d�>`�.��p�@�*2�HM�I45�䵐�C�+}��� �Q����B*���Г��<K���ED��r�2�֖��ȵe�s)I�t���Oi+��i����;5��./����@�޹.F��R��2Z=��h�	�ez�A���{��5\�݌��)&�l21��g���e	N�ϻ	�1W�fV���Ë8RJmz�D�_���K�%�Q��4�9�4�VF�y��rnD�b��	�z�αK�͏��<��t$�e�[�`�Q0�B����d*�^����>J�KhT�.��(�����y��9Y�{6H(M)��c�saO�H8<߾-���XeŰ�?b^Z�=!�Cg��5	W�_�#}�2�+El)�#+V����8��L������t1_��J��'O-R�
c*_:!��9�8$��̏�/p�H�#�H>2�M����>W��Ҭ������E�c2!trS��	���+�6���|w�s���]����J�|�b�mݓ��νi�س������}`x�/)ݙ�g�.��1A�NXŧUW��!6���O������ o�9E��S~���↩��4��QD�����c��o|Hg�@5���dk�8d5����$�s�Rq�T�Ҫl��q<���߾��|���܀om\V�ᩪaӓ����l�����:\Z&�!���M��)f�v�W�BBj!�֤�2.������u^	XV����ۏ�X�զ���$��	=9u��M8��k��&�����t�V�CE����	b�XG�<��@���G�^J~[�?�W����U���`�����S¨*�����,<|V�`�:�l �>��J=����܎I�ߚ�؞�E+��j_�9��=}�	����--�_y�(<D0|�"+�U�y��\jQ�����;M���ev���,���Vr?�;�o�%��NԪ\g��Q}��`':�����������;!�Y�o�/[^ ���Z$u��Bzyx�B���D�c�!^��y�V�ƿK�>�a�5`�?Kx�TV�3Z�΁�G�9��;KCf���z�X���z���F��T����x����w��m���FǶ��7wm;�ڠ�<p��k�[����y�>�S*��?��%��-wl�b�װ�U&��,�O�783�e�q�%FO�+?��Aq>�rR0r�"�O�ų!;��+���7L�c�^��pdr��!O5KL����f�w+��z���S��Q�Y�W��%q�dib�Y���V����Qf�5qy$�紲1�w�m�6yD�����(MfV��!<j(��m�ӂ��ON*)U���(����K=�{�%R�X22��6aY_�H\�5!
2�{�E������t�rH�����;�q���Ӟ�?$�0j��"�%Ps�R/�8�����lDb�1�BQs�=i���|�E$<Y�\��'�pBĘ���%�c����-�����>�N�®����̒��<<M\ʈ1�1�h-\~��c�P�L!!�z&�`�yw�|���U�:�\�!�T�!L�c���45�3<�
;��yCǴ�Z�Kr[��'"�0��5z�B�-G�j��s(��`�
�����ɏ���su�H�H�.�����j�Ĭ�R��hUl��G�d�WU���.�d��L�G{�?L��n��ۻ��%�]����li�q�kU���d`_����֕�f�����ި�����~�ǩ�΃��mG\0������ "�m�R@��H�����	A,�;R��i"-`^���!>���">�D�Sn�}LT�R�k�Z��V*lcJ4�\�D���9�>�2�^Hz@;��09F�E'ߢX�+�b���w�X��'"M(B+���Wx�	�D��L���TQ�	��5�����6�+��0X\'R{108��'~��,0X���#]��H���z�ѝ�����d��"�|���!M.��=��T�+@�)�{oc*.�0���q��ΪH�v��b��ōq+���S�J��fЌh��6w�0��+-���9��h�<�wl���|.�l��!ت0㔯�m�J���${�JN�Z�@ou��Y�;���
 �7�B�A���uu��>XaiVӕҪ���n����fL�N��.N�����5>rqZ��~��]��V��k{#�nR���a�溴"P��8���z��7$�y5�O!@å-Cu.A������rP2�,����-(�z���h� �Vpko���������2�\a�@�o>5=��X�_9��4��jǷZ�����T�i��řx�;~�I�R4�^�c�S���^=
\Q�ވyk�g0�����ݱ�9SjV�RE�ʒ$�����^�_tkE����'V�tJ�g�v�μ�PE�4Tu� ����:���Z��"�ӼG�����S%�*���C�^�ɬ���g�*c�]sN����Tf/(��˓a�����uxy�'%] pKj�j�P��O��?�a�ϛ�g���qXa�e��f1)��{&_u�}���Zk���t�3���u,���K�:z.k��#i�6a> F#����>;�p����d(�D̄=��}3���uJ�h�k�r����c_�Z�b��4��L`�R�#쮚#��J_(�i�"�59��d}
����:��n�zi,��L�̓��9wz�#�����GS8X�vG�Ǻ\_k���I�(;��%�ܓ ��w�����]���ޘ7���4�q�lM�`���U{�:Jv``aO7bI����y$p�wl�$"�7�[y�E�F�p���ii��S�4"�h��K���C�4���I��py�/�`Ps���1���+��{�ƺ	���
��-����* �ɒ�Z��7Q����K�O+�1}W��C���8�W���_Ϋ���v�8�<�*�P��W���.���I��T����Yу�V��B�m�u�D/J�ӶAL�o���a�D��=�C-�X�4����#;�(�G��,��3F�/�_��!�w��Õ��
Zt�E�# �cz��o<�,Y������"B(�,u6VB�"��M�9���������3�S��oX5�3�2�����-�~�W��-��Lq���������N��
o�+eu�G��7�?��L_+�s`#��h���NTQT��`�ONι-.����3d�_�<�rw�Ig���ۈ��[�j>I/���)#�6�	'�>�a�([�7���LÆ77T]̈́�~��U7-� ���O��sY����7��=:�%B��Q��h���%Q��hQ��.��5�ѻ�-!Z�D�eљ1���wݿ�ֽ�_��u�~^���y�9e��x~Ww�h8湟�jZL��
nH��	3��9�Yô7Q�I�8�g\��=�MV ��J�T$9D�~��t��Izs6qya9�)���]�7��䋥���� �����U�rb��)4[�K��#����IO��Fs1�1�w�(�Vl�w�A�K>�9������s������/S2*rR���j[���ˌ�U� �������m��?�$��B��vg�y~,6��9�A��!�d������*_���z�~�L���!�j��*z6�@����{{�#
��c��{Q8֙�{Kҷ4��rK�T#����	�����3����N��ܚ#g��,0%+�^v���?J�j�^��l���|�2�x���_S2���}�J	r��{á��o?E���~����ۡ�"h�R�ŕ��^����ϯ���=�EO{�}��< �y]���)��Ł��є!se��3s���'e6G��u�#+��?����!DD�f�m��ϭ�SGǳo��v�
D|m+�|�:��������GyoԌZ)��濋C�d���W.V���0���~m�T{q�y���{ka�㜜`�2�t�ǳh�M���gXJ݂�j���������4{�eՅt�����M�K�{�o�Ia2+��*HX���`*Q�����܏Gq��g�DP����y��������/C;����<J�����q ��Y����S��ړ��nT�����~/�rB ��QY=�tM��Y�ƀw�>dc=��Ǟ���\f�����/W�'G�g\$����EP�zpH7�0�p�y�l[�/���}>@�v��)�w,�v#�49�dw���Y�cއ�A����;�j�i�\�]��)���-=ݦ��c�3'�:�W:�wd�5=��Y9f����é���b�������D����P�ގ�r%����������)���fⰬ�J��(o2���\����F��!�5���	���ü���� �%�'M�_������ V~vc'X�ɒ�k�Iy�ʾ��'.ޖ=<D#�0�0��w�%�9�e�LK×9
����x��ѐ��`�ƞ/)���ѹ3��M�j�]i�.X5嘕ڴ�0?��V�3�(���ܥ��%���p�Hr�9lS��y�%�oe����D���=?!�׬a��),d� ,�$H��٨��U&�)���<��(�G�U����X���r;�P])�.2�>-����wd��h�[�I�Q�ɬ\�[��t��<����e~��)
�O���N��e���{��#��i~�q���O�z>�)��֒
qz��a�t���'|��He�D��mWW��e�j+���nxR�x>%�3a�Q�V�<�Z��?�����m$��ԍf��=��Z*�5�<��H��aYl�?O��|a�C��Tr��8`{f�Z��ghOo��}��"����c|;f'j+��;�A��Q�ܴ�F��^�(�G&���WAr�y���t�.��'�R��Q
�@���X9.p[u^�ԙ�z��'/����hB�@��7�k�ծF�XY����tL���F}�/�2��ת��3�Q0�M�.��w�:���)JI��tK��v�a���������I�ӆ?'�2��67��JW4�}��ۧ3r�FU+�'�D/J��g=�������=2��)=����/�eދ~&d/\�y�N�6����{�yP��^�b<�<�ciu��#t"�JRGI���{߆�^�N.	r:��Z�K*����s�Y�@�vf���)�!,���y���Z�l�@���p����ω�͉�
��f)���@�;�x	����B$�f|�j��5��L��:d��T�-��5�V|��wOM���hn
U+c��_V��f��(O��z��� F0r��#����)	��(u��� -��=j$�]±<߼�~(9��^��&E�o�%|3T�P���"Ku}��@��mi���`��]�~6|"'r:ȴx��+~�Y�^��)R3�F�� �]Cz�1A&Z֭�Q�g�`�=����Ee<���X6�D�����{i���ܠ��
���B�5��Q&��z���2�d�C��Y��d�?�6���Ҷ�QA�ƞ(�=/t}��8 ��T6#�8ߒz����Q���[Y��9��}��9a^J�t.�G�Q;W}���/�&�o;}.GX�[g�2�Syn���.?o@H���7\z��z���7�����b=��(��ȡ>
�u�-�i#+�\}�vZ��R0WY�5��D�T%�׾�2ݑ+`s1l���
�q� 
��N�=b�羫� (�=�HTD�|���(1��X�˶؈K*����gĖG�m���*Jˋ�_��D����q�h2i�6t,�ΪLi�v>y(�Gxl��X�V�&:r�ֽ�ex���Tj�a�51�aY���2{P���aqC��6�;q!\����8�~�C��м��HwlC�2����z�aҽs����`�%�y	P�2x��ª288�U�V��+ˀW?�:z��d5j�[��&�݉3�O���[�Q�#x�Y�v�^��+�ؽ�� ��F���L��h�4/��Q�R�2e�l��7��{:�#�#/�d����%��6�\���D�����2�"��?*�^��QNf�:ݗ�ۜV�b0��o�yۀ����'*�k�|��G��V�}��ux��I���)%]gO�N���9|���;�#�z��"��8vjț��p�����
���ahǂ��=�;IQ�����%�ш>�M�g�[Kα�Q����:�R�~�aQʺ���e	�q_����\4;dAH-� �g���:}:�fSd(�'I�+o�u���;'K��(69�ԦLN�J!��,,�_p,]n6M�a!;�Nl��Ǹ�ǃ����]&����C�y���wAGy=�b�����0vz�8�&D�M����CG�o���P!ú̾�{h��6�JɆ֓1 �=3�{�kC1걸1@X�WvC��Yo��5y��b�2%�c�Z��Q�=;�Y4�UY;",S���J����sAK�T��m�-�f���y�� �$����HhBl\b���@S�Й�8Tɮo�v�ˊ�!�F2�ͪ8�rԕ
�Mй���
�縭�����gr�zZ4kL-UªJGv9����I���Q*}��\2pS����� �@���"ӊ*���Aj�o��ΰf�^��˔��)��ܡE̯�>�\X��\���^�FO`��*zߞ�1�����G����2=�Fo|U-������X����f�'Z�Μ��y�{��9���v�"�����o�B��i�2��?i��h29,9;�������r=�m;3ѷB2�Ӫm��T��ܥM���K���l��+�>�/�z��%.��`�?W�$hXoy��ߕK
D�	*�����-��\a�{�)�M#<�;C�n�fP�\���Gs��0Z����T�p���Hp�)�dS�Z�ƭ��Ρs�S����f��ٍl�g�����$.��(�-�ؖC�m>����V��c�4��&�Qh�j�:�4�0���Y�0��~�������,iJ��J��q�Q����|cߡ�@_O���~����Z�Xǝ����1��z�BĢ�����������Zص��[9�/19�+:\CZQ'�z��g�p"66^g��!��x5����R�,=�g���FWMzZ?��8�!fV�gF�bz������+h��%�:;iW���?��Rƅ|~Ai�wQ\��?�/���x� �-u�N�X�|92�������-:2�O�p�G�]_��L/�H^N����+��Ž+W���8xvz
3.6���E©!�#}qm3�3�OQ�j���*j� �y9������X�9�q�����l�����Q�T*m%�T�rfw�����b ����B?���F��=t���IJp:q	?��w��H�̊)r�U�����]��zX�c(I��Q��U�H��������	2V��K�q�r02�/�c�	�~{
a�*���=w)�#�9�����h*�=@�;��	�'!x��:m[�ڙTd��R�}L����X��uV�駐Q�����F��'L�v���e�ڜ�u��4���d]%���P���4�D����|;h�V�R�4���D搕g��Iο��ճ�1Gq+��I�ȐC��+نI>9v�a�߅d8�%H5�>8�x6&��CNU��<I�F�h�.+�Yf���%%�b&i�D��!���V�켿�"Z��kE�#�|EY*t�t)?���<�Q9�Tb�]�1�2v����i��&���!X�Oki�QR��|鲰}��ǟqho���L��q�����S��;E����7a�K]*Ǵ:����2�!*W%K�u�🷉�c"�SdH�J�Df�^���bJ��	��B��g;'nR�X.�qԋ>B��{u�F2�?V8vߺ�Ԝi�T���PG�=��ݷ������?���'Kl,=n�2u��s55�ڰ�mqK�h�yIl�҆,}�-�h��1L9��v	/�����ތJ�+G�+�ǩ�'����Poγ�>�eb������ s-Z�Y�U�'�P`k�q�T��Q�;����%�z��㱎�'׋pvC��'��5�*N�e@�x�漬X������I���cs����Q�	J:�f�g�[����.���n=.����T��!+1s�F�((GG����Sy���AyҼ
���*˷�[`�Sf����fX��ǔh=)�m.@y�z*�|�śR��}a]����hZ"D�	�@��A!������G(D(��?ģo���uU��~��@���::b��7!w�p�u�������6��:]i�'P҂!�̸0D�D�=��ga�+�fB�3pK�y��d��OJ��g�%���c˓=9�8p��8Z���D�A�O��Ú��~�+!0s���7,��~�H��&�}���A������7=1��
.�.MIs	�]�������ۯ����O佊 T�Dr��\�{� � 0tg��ȃg�;� �ms�I!�_�G8�k���x'�[W�z�+a�2
z慈�e��2����W�#���R���3��c�:O͈I]ԍ���څ�T���a����g�cb�T6�|��KV���uլŮ.GLiON��k��j3I%QA�m�k�<9�����TA[�U��DY�sn�:��V #U�~�f�<_��� <������)��9���,S�p�r=V�hEʿ��cm�[�md�n�M4����1�ٟ�䥟���T�Ax+o��! �d���Go�p��+���J__��G��A��ȏ7�̳�*�C%�q��(������u訂����WU����2G1�2� Δ�v�/5�����	0�MQ��s u�fy8��vr�����!�ND8�BN����LL!�ce�0�y���\64,`�}�Ɏ_��qk|_��6b��ě�e_��E�2;n����E�Zx��t��J6B2��{�/y��a���IGɸ�� �rN`A�UK
��x�����u���F"��OT,?�_�Z��|P�OnH��)U%Xz�o$a	�����?iʀ�K��,��(qe
��=L.v�v��r�J�����z��ss�f��׉�EG�-��K9p�ɕ�|��n�RAy�*l�W$�}�,�x�����'�)�� h�R�6�(�H;�ӭ<ͩ�Q��j� �n�1(M�혅�[��[�_o`��Tu�q�^0
���D&7t�T{��������]�r��_�s���D���BU�[�h)^H���)7:�;00J�G�^Ҝ;�ۑ��-o� #�U��%7�G�A��x/�#�**:�!����X2ӥ�G�f�!������qP�x�1lw��2W�̲�Ih��pX��}��klodw��^���E�M�H�������u��PH�����ߊ�K�����#�+C�r��2��p�85pe���
;AŌJ��(���F�^��ŭoJȼ�V���~|6�=a�.v��`D���H����K'�����Vl�Y-�	+ʪ��ꍉ���@�Cj�^�M-܏l�DO��v�=�������qӒ�����J�G���ĭ����l6�	$��3g�Ǒ���ts#����Ȋ�$g����f�C�<�[@D>)C�U���\7��T�>�0�jv"���A��2��s+pɗ����i%���,��+'IO�hX�*i-M��$�&�0l`�"E�$i��gz�2�����y����އU��^�(��v�&r�i�}�g�U��РL�!�<���
ua7W}�E6�da�����&7Y�*�-<�wU��ze��c��g�[q���pR����77�FQ7Q�^�J�l�
 �9+�V*����c�[��4�߶2���o]
Ͼ�w�b�?K<�E`�3'�\W���ڔڗ�� �*@Y0���"	���:�✾k9�̜�U��(�.��dLF(EL�l�K��}'�:D�{p$����R�tQ+n�������P�K�M��e��מ�6ss���Ӕ\%����A�K��JD`)�{Gj |�G���<�������oW�	e���r��Pª`�\�����yv���=��F�+ɪ|�#�u�T�;�}"M�����x6��w�ٮ7��,m�l�n�WD��0��J��â��}4��w� ��R�O�3�s�Ӳ��t��3V�7}ecN�~�]s�#3��#9�ȒR2��o�]aĞ��h4Ů��B2塵:����{� A��/���O��5�F�@C���UyJП�i ͛EiU��tu�?_F���:8�5F�H|�S$F��68�����t�r�-�N����e6���#������w P�����o�j7�c|~aƭ��p�;�%��Z�J��u4�s4��Y\����W����N>�u(��g�4M�����-�\-k�df�2Vf�b�y�5r��+#$}�Zd��}{ ���1>.�N`y��̝^a���]��cU�$��G��K~ƫ?N��S��>�E��/�p(o�M���;$6f��3�>��0N��;�;��a?41[QJ��6|0ÙLT����W�J4��L�c������AL�f�ȍM��;�yXk�El#.r�����U��|~S��=���pJJU�����=W�_��J�!9�� ~�� ��61,e�ҡ�B��t�=�S>�tm	ޡ�j���)[w�����qzT�t�+���cj���vI��V�̿�Մr�g��\��>�K�ɛTO>�Z�y�D����	�4��� v���cfF'ŀ=�{]�P}E�+o}���W��VR�D�����yo��Zr�ݕ%瑅k�����g"g�T.L8�)�!����	AJ�^�05��U����c䦥@�>n ��P;>��{@Hw+��61�%x7p�$�ܧ���F7_Bw����#��e�j��2�x�X���w����"� ��_��Q=ֱ���Y�˝���m�����;�:v�I��;�*�
x`J�N��䚿�@�Y��8��C��r[��7V�n0	����a����_��8��&�Zq��(ʸOA�ׯZ>$9�nȴ;CM��� ����-��<��o��I�5��]�n_o6���!��y#\�BB~�1g�H�^3��#��U�[vt�ҽ�6t�0�NAP�� Q�j��k T{�k�-[N=�����I`���GN��*��Z!qlو��P�����m�Ŧu��[d%�CC����B tG�A�m��a^O�+%ĂS䖖?����Bd9���{�j�����Y����jL7h���}w2����ɭ�^������/�\�g���|�dq���[�$��8�cf�����T���.
:�����}]��nG�9�܁�`�,�{1����?e]�$b�E��k=�R���&�����v���ڤ<��z@����,
��Y��y��i�v���I�����S���og&(��^�#>�>��o͂�Y�U��Μ��8���?��3H�~�׳ޫ�[1A4₮��2]BW�;�&�V�I���-�}=p��({�ޣ��v����lX��꟏�P��ˌ��2&�V�h���,�� �&���>츎iz�q������
N��J��V��k���e���2�>(������9��*p�-�	Q�g�)!��Ufz"���X��B�>�g5���bHS���xJh6���d��
Nctƕ�i���ҟI���	�nUh;|��[O���>Ǟ�6���̤͍��`-j�37�sw��JT�G�m�i�������:Ȑ��e�t1:�X3���$�������|=�ϧ�9L���C����=A�K�cZ᷉ur8��O�/��ZG.��r�n1zMQ��&	ñ}Qy�'l�Z�9[�?�C\E=�nǉ����7����8��/.o��O� l�; �O��rK|K��"o?L�uB�~A�k� ��F��-K�%N�k�D�(x���D^�}��o�)�>Ѕ��8%�Lpdʚ�)��uS3���hP٢G�8�g��u�6�D�S���̬��e�m�?>m�`t�R&I��3�b��Y�'k��6��qdz2a*�@��ȑH3�3��$
l$8>���x�� �&@�(�r��]�I������ִa+.��'&*�j���
��A2=!��g��I��f��(J��bD��K�A_�����;�%s5 'c�Oǻx�^ARe�_{���D��Q+��k�/���>1�B�@����C�����3����2�%���P��#N9б����^�ɩ%��G�N������n�#C�G�w��Z�a��tG�R[��_��4��J�Nd�?���Ƈ���t"ΩH��������⋼�HE���g�v'�����q|Y�m����I8c*Q$:�o+־��N�Ǌe����Cy�"�Ś��C�k���l:g��w����;�g7�)��M�~���I�K��; 	>���O�����i�bѤ��E#�|Y�q��r��AC�:3��;�/D�΂�Sz�����N)��i	s�	�q@n��@�wQ��ְ�uee��Rը���iV�UϤ�7F ����Tդ�gGߖkT�'j�ʱ���	�ػ�/�av#��K[u C�SQ@� ���J��C�O&iL������SF�N�|�&��O�д���7�������}`���MO@�����4씄�����k@S�"&�Iak1N����a��c�?�D�盏7�C5�˹��{fh�.�,5�j$�gu6I��c����)١N��T�\��t��_l�M��,h�y����g�N8������K�<S7��>��
��鄙#�7=�7'#��}Gz:g��(�=�WG����)HTީ�+c4م[��̸PKmO�M���`Oza�a���\�YK��ל�
��4�V���X��8�]NW>{Pj�	f��)$<-]8�b��
ܛ�����~ZGt��R>�`���Ӓ�F��6��W:fH��/w �۞�3dIO�}�������<�S$�3�K���k|j���	��G:����r�M���U�0ϥV����ܐơc�QU3p�~�KD�!���Y��s���B~�4�	����ed�xSW�Z�4>i%8��������ĚZ>'�1<؇��I�'���!�rL;Rjj̚���V�
��$��F�%��x^\�|jñV�=u�YZ�%�C���P�$��:�8���J+Yg�=�fv��iOཤ��/_6P���Uؗ*4y�p$P_��N���-ɰ��x�E_���:|��h��W&һ�`���Q�]3S���H��*y~���0.��b[J����݌����[O���	�@��s�ɑ��;�R�F2�$tv1h�ٓw*������Kؖ����O���nǯ���(��WN�mT��7%Òon�pϰg��	W��G�fJٳ��40��h"��3L7�f���U׍�a�/�N����f��(��{�?0P᷆;O��m��z���w =�B�4�~e?S�&!�}��u7d��UZH�ra.]`A\0a9���7�.�E��H�.�Х�7$�/	����(��D�z(ӳs�rCy�Յ)�y!�a���H�J�!���}8s���I8������٨�O�J�P׼���z`��
���J/��Z���\��'��L��1��\�vg�G��	�r�<ƴ�� �5�K�d:��*q[ާ,���z|�Us���{�.�ƶ����/f�j&A	W}d��!)���`s�`�I����6���� 0��;(-�ov:Ls&�³98A��@�_��?���v���H�֭eL�~�"�of��u+��N�2��,�F��|Ur�(�IYJ;J=d�^W��v3�N� g0�J��:��`s��{��������.�<�l���&�Q�P��ŸT��4P��z�|��m���#����n[C�H���qI��=G����*�֙Ӟ��G6�g*����̈O�����oѲ1�r�0���dK����J�w!��`D+��?��f#Zm��q>v���fB����~���W������^�2�-ըM� ��j����*��/�6��ŷRg�>L��ٕ�������nN?��`2�X�q��5��Q����zLm�L�Ԝk�󚪰��[u�~C��_w���F�N�Y*���v�T58'2w�F�X[W���qqsh�Z�|k�'=;︵��#Kz�jĨ_�o�I�BP�r���|%����_U�ם�ق(j0tB��6��t,�����;4�R`��p�z�ь�Rn9��#�P�M�\���f�+�s{n�ظ�z߿<i �ǣ��H7��(�PQ�,Z�qh�����d���n{ݯA�Hޕɀ␾a�Fs@,6��g�@�����(�����&�}���QAղ�����԰"�i}�yp�=�� VPF[�H������eJU��*������_����Tu�f��E��?����W�W�ro��ڸC�LMZͥ����LH�w�y�,o�Iѐ'M�ɛ,�/�繸���h6�K?��Z���|�m��ZK�N�O�kV�R9ӺnY�ƾ�YY(�A]U�Ĺ;�����L��~��zj�F;S~��9��O,Bx�8��}�1x�[T!��a���� ��>�v�� ��P׆5��\���-uVa�����惉C�6A�ݖ	-�� ��h
�%C,g$r���pټ�r��E�1C��=�+���\�$������{�����\�:_�i
^��.�����&JF�/���2���H	5a��%3LW/p&���.�]NH��ϳ�E2��Ӵ�Y�3�"�?�.��v��������,��H-�XO�Y?�ll(`�u�f3���� \�e�+X����yr����!w9\=��m�zkՄe��,�.�@�^K�k�~Q�bJG"զu�h0��M�>�az����"�����Ǥ�]]��rZ�İ&�^�*GK�]���C����������sv�
V��iF:�|N��o�P&X-�9\�pD�Jl-��mΉ���Y���Uy���9�r⭄��4��:�����i�W`�SO&���N���_���q�����.�Ǉ�?�^��|�eŜO7x��޾��jg�����I� �0�p��D/p�M�i�(Y���z�I�%�M����Ǫ�Uu�gh���Awߺ���i)���s����v�)��{�1�ܫ��ll��&���_�g��x<��v2J[Ϛ�tvmz��t���˯g5��7Ҹh�;@f��!DLă���z���p��{��ceO��Y)�FUқ�á;�gf���T0���.�W�:� ��]����UDMY���a�'g|��0���2Y�STx�I�h�K�S�X�8ߊAg�łMu_��k��Ё��ױ�-�G���u��}4�ڏ^|���,��%��I�|A�%�w���^KcS�������F9��%�oD$��D/;AoNlxpp���ۢW�z�|�rlT\�8�+���C����4���5k�+@�iar�8�;���6���ϟa��&��EwI�[2��fb��Ҽ������� �$�����la-��!���e����.r	��7�����I�iP��,l&�XVs�I�t��^��x�&�%<M!�W��Q���*`�T��I�[o�=�ŅPE�W��� 䣊x�m����-%�P�β� �E�J���M�-�� 6~��8�*�3�:Ȯ�4�.$Q���+�^���7${p�9�8�"r����&6m�� ��Jh�ȞQ�{���R�%���Wᙛ��Ԡ7���h���]�s����Ҿ+�$��c��,/f���ɳޙ(0P`���p���S�-ա� M_���4)��*�y��V�8��S�J�V�n�}�'S��Z
�/���WF;��t-{FR����Bj�Zm3�a�L�L�&��&�\�I�_w����[ƕB�
�S5�9��< ���Q��W������^ G��_g?L�R���[���p�Q�H���e�@��:e'����
�G��1�r�Uτn=��n˧��^ǩP�/%5^�g9�*��)d�yv�+����JXVZ�];��_q���K?����K��UW��������y���L�w {��VބN-�raT��[%��*�X��H�t-�(�&C9�a�L�z֏kA,�qH\�˥ܛvOr.��.����ޜ�)�0�~��5ظm�>�{�eB�XI��gSaWM^E��[&R�3����,.�����kz�����sj��'�3�?���x�3���/�DQ�&�w���.�𐢩#{XQ}z|C�gD�Ӂ����d��,��
��EP��K7P�2�E%��3�1�1'E�;��n��!+�����9*�$5"��5�����y��q�m[�xl��t�[Mj�LY�}r
D`Gp~^z��0�,��}��-o1xnRŻ.����l@�m;��U�b9�p�!�}qpv�+	H�'��	��̳�L4Vr�S�Gѯ��YR��8?K����
����5���	%���<(ߗ�vо�Xdr�G�,��2���v�x?����3tC ��oTb@ @0���ᱟ�S����_"6�ߊ1I��.6=VM0$�TP3k��kē�����`�TF�1_�$B�~N�c囀b��@fy�dy�kEՄ�I���F��c�~{M��'>�R�wn|f���1=M-�5ɍK�K�?~%BV���W6�]�j��fMؒ����mԌہ�Y�	T�+���JT�NQ�P�"H|m������.ϤB�F%&�'T���>7����]�iނ8��-�i�S6&V�-��{�xm�A���R���۔^��a�����.bL:�l�d��\'��*(n�ϊ`ճ�SC���%!�i�n`�gT�s���z�締�oq��2/D����y+#�25@��tF>���,v�)5�!��13L��G`�0X3���������ZP��(��t��f�z�xK�xZ�6Y0�P(���5.��'�~�w����Ѯw�̢k$��-�a�6+,9�s�H�|g���?)X\��62H�f9GP��ԥz;P�bk�w8��"9���x�X��&	�r�W�w��bht��l�1�k&���[��S���c���s7�_�2�0�&�������ƴ��pA�$�5|?�{!�_��o����7S�X2���c�}�L�8n�+�������9�/�����x�	���!y�5�{*��bG߲�]�o	wW���ʻ@ftN>T�o�υ^0����+�X��� �Ĭ�m�}��K%쒙>��x*k4x�;�V}�+�B�{1�7xX樭��K��6G����?��߾���� E @��i��
w�LZrTkK��ʉ�k����������7�x���LDn��*�Q0����L?�&;xf�~���Wk�����;����`�Ӄ�.�@Fr���)��ցA��_���"���������Nnz��>j�E���)	^�Łf��\�J�ө�M�`��ހ�y���l�������X����ϟ�)��|��jk��q9L8�bi@��������C*�K�o?VcY��/����w��y�4���N��t��u/�#B���!�/�41�5���kp��F�d��s}	̷o� I���F�͜���/�g2��C���k9<������5�.�!x7ˠZs��8��=oӸ"���+Pi�|�G�lRbZ&C����Ա��X���l���_����N��������=T1�N��5��z3f��%�[�x�K�A[`�������L����ܭ��ˑ�h��b��2��!<�K���z�"�����pSMBm��b��c�'�J^_�;��gq��7�����}W��\ex�����)�]����@��;��eK���2`���Oˉ.��n���R�|<_N���(7���}H�c���M����[���W{�W17=�w �!��Pd;(��`g�b�T������{��q�H��2�?�vw9cc�؃��qu��v��S��x`��bL@�11}���� �U��<���tf��`�1����o0#�����T^�/�Fi���	�l����BHЃ?���,����s�tz7�:��&�)I��w"t�@��vH}q���'��c��{!*�����S�U`���I-#9��|�?s��I�a��ٗ�0`��R�t�愬�6�gLL�w~2w�rȭ����U�wpr(�ܼ�����\A��C�v�M�����~k�sΞ$c��c��0��{�AH��(h����blT �Ӈ2+��1I�ƜhC׫s*<ğ>T)tg�#u�˲�_~��e���2��H}9���e���rp�Q����31�;4�Q��^��V�68�����E���+m��x[�� -����K����.��$L�� pl���@��.�^���j����Ub6���ӿ�����G�ҿ���� ���j�D�Ӏg	����K��;��b�+�;iS�w ��)�QzJ>u���_�0v�)�� i�1�$U�
=D��( �}�Ƒ�!T[�|����3��d�?࿼�k���_p���_�?���������p�������/PK   s�eWV(j�Y lw /   images/89e20355-1f0c-41de-86ac-b21eed32d9ff.jpgԻwPS_�6�)UT�@�z�����[h"�ZT��Kh�{K���Q�t!�J���TE�����|���9���|מ��g�{e�}����_�.nk�k���� ����
�S-�� �� �  � 1� ��3����b���O���=��� ���ޮ���� ��H�KD��Eo�g���b��s���?{��� �HH�HI��H����nRܦ��u��-������c``f�fgf�20<|����/���.$*�'������"rrr��w)(��130�����=��&�c�-b":�:"b:��� �?�$%"�� �ALBJNt�V�6�����)�R"�떀j���<S&��a�pO���KzN�g%�&�$Tn��ݗ4q�L�6�rm���迎@�	2��JQ�k{�	"���Tґ<�#ơLzW��<�_���i%\*�� T��=�� J��D��1���+�����@��?x�����$$$���៱��IHn<Ҿx���t`�O���7/�w�����?_O'���4�V�՞��
չ�?�/n�ik�����7ۗ��ݫ��Y'���_J,�����276��<�/v���0�����C��/�H:�5=)�^6�	s�eV�o`����q�o-�t��E|��޾�Ɨ���I�B�}��A�F2��_�o��x���9!i��%ZV 2���i�ךk|�����eTQ���U���jه�+Mt�Po��}ZbU���� �'D�������n��I��)�߽�Bz�g�"�F����A'g��J��iӌ���!W�G��t^�=h�s3��+
թ���H�3��H�5=��ڪT�?��t�������Ey���d7)�����?���4fRx���53����qzZ��p~�Q�����c	���t����z��ƫ�	9��x7�-�aV�y�Nr4�NH��N�G���:Uq�8�i�7�ƛ�|R���Y#�Fbz׸�����[T,����H:q]nf�&QL��9&�85ds�M��ޫϱ!q��X�/��"�u��1 �9E���nb¡�\�>o��6лo���X@C�*+�:���A��Y�f++J�Pe��m.����[���eJ|H�PK��x[��84�F�U�XS6&,�|f9��v��*n%RU'��9fԷ+H^EUx���_����Ěe��n�l��=۵a����*�L�Ѯ|`��rI��m��Cª��Q��7�$�v��֯Eki	�n8��h��.�}h����ngC1�懛�(��Ň:����q�qm��O}ʕ:��OZ�� i[Q?��ir�
�`����ZK77��E�'�UC6}���.G��\��r�5�J'R��Ʃ9�lǙ���)&�FN��o;7~Iݽr�����_W3|�m�l�$�Q�X��28`�9jf$��_�*$Io{�����8[e��9��yf�(Q�LhTff��ߒ�=�=�{��cDq�B9��
H=�c�������
Hh[q��<�̲�[���vG����L	���B��Wrk����~=!��ۅ�I�� ͽHH���Daȃ�e?mn��{sL��������,��T��/�~�/�vع�ؿ )_�k�aR���j����<$�B8��/�S��s�Sf"i�PX�t)�h�\�JxF��0����ޢ����:�v�bB{;݊J(�%����Խ�Xcm
��rM�"�>븚���k�坘\� �F�#qa�[[U�^2:�=�1v��̩܄�@���ߛџot(�oܞ,��҆�?Kr��=�*��&|a͒e~}C�u�s��"3ϺT��K��C�-�r�$���1?Egj��}�����=�m%�Sz��#]ujq9O�O�2�*X���ƽ9�\{qD��GH�Pj�IU�
~1H\W@Ê>w����T/�:lop��s��0iY>0s��T�0˿�R�y��~Ûe�e�"���l[e]�����j��������²�I[�2i�B)����'B&�����>�w�v�aQW4䪱�'_�G���x���TQ��(z���.,V�!g��T��"�(�S��ǥ!��N�[�� [��t+�t-+��>��ꐚ&3F�1m[q[T��gt��Lǡ��odY�^2|5��LWu�NcB,<ܬ.t'�ӯ����89����nWn�*]2|&�pW�b`��1��!��歃[v^6w��	�	��	��M��ڜ�l�i�y=?�y�O�ux�@�����U�Hƶ[��3��J�%U����x���W�>c�tmV�����bI/�Y�:��1�c>>�VS�ʊT	����Dy�E(~=8)�;D�<,��3h�V&�����$+f��¦�S�}6gG{Խ\��\b2���Cs{��LE��RZ9�]8��J{n�D4}�]u,=�F��`l���k��:F_M+VMV?�w������@��3`j��?�udtۢ��q�۷Z���w���j�I�(�O������?��
�I��=�Wȅj.-d�C%��x#�_4�\ۃ�с�f�Ш^�ʍ`�3���ɘ�B��l��E53x5��*���5aj�	CK�}l�\ۭ�_+>N�L�!�m�*wlQ����kz����A4$3�
��j�~���ހ����fx�8gx�"��y��tb)A��]���:���k"���r[ u�=�
�������ueg��,�����{��Έ�aܶ>u0��.x��R�ї�t�ͺ�&���r!�뾹K �f��d[���1e��Y��) -�	y t|��#1M�����6�d\�ݫ��Ū�֖\
�ٯJt���y,gt����@�Z;R!=$BiY�Rm�x���ap�q��Ma�5��%�S�cRN13
�WHz&W�P>�g ,����]B�6�gXC}Qu.u9M뒧C.d{����x�5�k:���B/ՙ���B<��f���y�l��\��3lr������U�C��u���ގIړ��˩F���WG{�Wp�H���<KG�J��(VMr}e`�W�90J�,o�k���%9����m�V㿖$37oCʱ�����T�b�n�cќi���=)�_�;B~��+�IˏQ���Mm�S产W���
�UP �i��Yw��9ȩqM��ך��攫G���p0vN�R\�����\����W���u�f��
�:�g}�d�����07�+���M7��u2�q��zi��\j'R�V^ݹ^�a���>7AAuI�) ş�l��U�4tͥ���ݩ�e ۇ�s`~zLU��-�І����#-&R^}��5��ݴ������@��=�&��sv�]����{�fr6�r6���Ӱ�6M�%�[ۅu\4?-åHĳ�Jz ��#�S�pRU�qU�_��K;J�ĸ���j�9%t��?�V�]�TL�IS7�uommLI��S�����X�uh�Zg؆<AV���[�ח�"[��nw/젥ҋ�6S��9�E��r�Z���2�}K��Q���죺<,9���td�I�
����ґkF޹��#�`F~���*��֏�\���k~�H|�\�[�۪C���V2�sk\��3�ˇ`�����GУk����\��em�ۑ%%�Y��	s~�4+;�Tk�XA5� ��QQ!�:�V����@W�<��b>���7D�l:	�E��^{l ���EZK�f �F�Çy�����w�-O��`.zh�C��4��X�A���05kf���a���	��6孭WS$��x��{�Q'����z�\��ff��Z��2ʸ�
��9q�=��1���<(���km�4�yGnOi���p���X@O-Tљ��e��0���Ȗ��F�s�����&�����뗋����	�Gt��.���7�gy[Q� �j��G�?������`oV��=�n[?.)���)�;ћ�zv�-���U�ٚ��=���*�.�5,�#��K~���0K��U$.|�j�s���Z}�ӧ=���F���w��^zY����o�+�=�.25�����#
Jt~i��6�_T�N�|�)c�ڈEe�%�
����hX�A��P��U�%z������Dޖ��Y��8�u`��L&fM��R>x�Ĉ8���_]Uꨟ�R9�a�㍮��"�Z:����Q���I���A��R���6am^�[���S3��a͎��)��m�#��NAU|X��xj&��9��4�{�:��gQWZ���-��@��Z]����&��
xݕKk���h|�p����Kw#SߊVa=����x��"�GM��� �0d�gZ2�Z����RPrJL�������gv��(9[KҐ��\�����l�D�Jҁ��V��p�SR1��=G�S��pˍq�Z��`{z���[��J�ހR��oَw'�}��P�h�L�D<ک��E7�<Td#��Wm�7�����'��Z���>�c6�����*�Ǘ�x�)��	���B�4�����yJ�='d�C6�{Yϟ@fOb��i6,�c�kq5%h���������O����&ua�X�e�{q_�f��
u�g�hhH�:v�*a�Z{���� �����э��-��3��P�qm�x���4s&��Rbln_V��$0a[�̏����R�JkaI�� �'kO(�F�;��$l��!y���lh��M�P��
���z�}0$:��G�0ʀ�D��G;���a*U
�Eo��%QЩ.��s��ԁr���oq]Hc7�:'�ۅ9�:v�/�9m
TJ��r�c��$Ck8�[���K*�3dv�&�����{�p�fv�M�d=hw�Y���3�4���� ��rZ7��rgF��U6��XhϪ}Ϝ�6��K���o�N2�JV5F��l�؆�VӜQ|U�T�eW>��\�oQ���~�a�����ճ�s+6I���k��2!�k��(E�1+���UH�?&�}�<���#�79�pfZ��Q>�.��#Z�cy̴�J��N��yf�d�9m�\�
�����R�r]Xϻ]:Խ����2Te[�\�\^w�\je��Y����.�#��o��Yiۃ[f�b�'�Y�:�/"տs���v��q0x�P�JZ�W$3��E�6�qPBR3�	�j��L����ܟo�T�t����� A���������Оl1�̶���,#Y&�$��eD��dW>�<u�U��$�O]�[�azd�,Y�@���}IyԲ��W�qx�����E�o��	�ۊM���>�3��ݬodԯ��ρ����T�|B�v��$ԖZ%��?����[�5��M�Fq\�]A`�O�D��"�Q.s8 �6������j=n�QN��wD�sf���ڬ�#�JAtsD��6�w�yѝ߃�@vym��=}%�B���X�,݌BK�G���d0<ɠ6�j���n]D���u����h��G�9s��);��������*A߰����!ɣ�PG��Ć}�LAw�B��H��2�V��& �G�����ǎk9�v�F]��)Pf�}o�j�n#9�⛂��д�"�<��/��f(�1��/@q��ņ����:�&�T�e@���6LƯ"1�04�^��3*C.��e��M�s�3	��`HxoK�.�J�g=c�X�ͅ��"����+�M @p�֥i}Ӊ��ڣְ�o�4˙ts z^�7��Lߑ�Vr	��/y
B�e��EkΟu�pt�g@P����V"(��T��
E ��0;��>���d�����G��9��|s���H�����X1q�ʔw:���S�x�'e����S�j�p���}1}���A�wE��SY��/h�-GFw3��%=�ȶiJ�%���t����ں����?ل�� ��Ǔ���\FB�6_�>�
�컚<�G��4�.Z���S���D�]x燣��DE�C�
�Ī!h��D��@m���l��~�F����n3!�wz��GE���荍�A��(���t� o���}O�� ���h�e
I]Q��Y�FZ�4��k�A��f�1����ʚ�e���7��Lo��8�uZ�L�����:�Z*���RB3F�Ʌw4�&�p��n�Z���k�>�*e�]Sk��ʫЯ5�Je�dWP��CWV?*��l��jr�ɛ�Q�Z�Y%S&���g�HBs�&Q����*�Ƙ�d)B���
Ԑ�WJ�x�iL�0��ǎ�Mx�h�6��m�ب5�@�.(�H���<����4�6��b�����m�'hm{L�lv�c�l���2ko�R23 �S%&���t ����WT�\$c�7M��\)rv��`[�j�������e���2oP�X�A�M� ��퓺�^�pg-�U����Y�o�ҷ!>�D~���)1�=�%�&O�����{������]mV��B���?�����q)qt�<������)�ḥa͍�S���Tt�TCY�[�t�z�]�X�������Z�G�l~x-k�$�a��.c!1C�\l�c�j�*� "�[U�����Y�J1a�E�T^��;��P(�1uu���Ii��c�	q�l����z��N�[Uw�x@���ee��Λsiev`�2�Q[*��,��u@6���I>=���؛�Q{[lti��g��X��k��;�b^6ag٥��[�0�9�T���O��~?�u���sJ:���xɻ,���[��y�tN�̒{�묑U9Bn���2��&wf��GדM�l��M�ނ�� ���ŗ�j��[b��6%�B��=�K��v�p�ys�GeӪ�۴��d�T>��L1E����.P!����h��_h�A��_�l�կ�)���X� ������`��ҁz*na�j�i|א�۟[F{�{��
'm��vCƦ�Z�jߞ�)��<�Z�n�W�|���L���*wcC�Y� &����z/�%4PsG9f��x��
v.B�}3P�9��@� ���e&x�m'��m{f��	��x�q9�yΣ7nP��*�_[Y�\}O�ǜ!�پ��
���ှN`D?��+���J�t�l���B;�呦E��[SF�/���j���`��|���ku|���}��i�I1Ձ�����L��7�X�|ܿĭ��#nH�׵��m�Z�#~ī���K0�&�M�[��ăX��?�4{0i�%�6f�J�@ބ��_����(87b B����f� M��[�E^�A�VB�R܊\���|�Ύ���&�������%GTq�/��g�aSҜ?E���ºVRo�e?m�&�n�T��ɀep0��|;�ޙ��Ֆ׈��$����_�66q�UWY�,!D�S���jԶd/A��8�gx���j[��S{���N��r�ܩP��E6��O� ��)tW�ě��X�q9*��V�G�����c��z���?k2����2�%R��V����`$����P��4S½��f���P�|X	�DK�[�Z{4 ok���hJ�>�Ut��������wSKP[���V��IIT�ҍ�v���D�ۅ�AI�H�IH�R�iYiy"D�:��S�169� ����L��}"�R�D�Se�
R������\GӤ"�Rc> o���]�` *��,(���tD�C�A�aS��?��_c$��&�D<Fn.�ӍƘ	սw�����}���@�Z�[iS��>o�"���"����S��
/��ܗ2/�H�9�Ip=�	���{u])�1�
����H�">uD~�Zc.,A�D�b�)�N����[�o�<���n<M����Y�ʂI�-;��5kp
�|��0>]��a!4����@\r���6���l�fs�4`�>G���YЬ��R}����mر����B�ؘ!#T�Σ��au�`��A�;�&�g���N����\2q
zܶV����p���R(�-�2�.u�����P�<�?����f׻Xȍ�N׫p;U�?�Q5��(h�B�W�e����%���0i�i���W|�<����N�Sˑ,��S=�И�����Gq���~԰҃2e��br�s7��*޳P����'���q�#v�*��H����|��e�bV�����M���#��w!�IãE����ao��e5�ឮ�o*�}����;�*<%5᷽�lg���'S�v�w?��L�ަ�b��6K�rjŵ�ͪV��6��x�-2#�r�9�6���Z��*P�4�Vt��KJ�INLZܛ�� ĝ\gg����K:%1tw}���|s�Ń{[����:$��u��>pK�Q���Z.�s+,9s��F4�I.�([4T�ޒ�nh�݈Ħ�*|kh�?���P��H�a>[���-��i*7 |�J�?y�����#�SΥ� �����sb�@�(�7��︡I����-�Î#�c>�ҹU��Q�U��X��u
f2i���\�8|��a%�C�����Ϗݝ{̊�c=���[�X��mc�[%1�>���N>�X�:�:���W�����1�"��lh\$mx�����K��L������1��ua�+�և�7�g�g���5��1�3
��-�_���h�y7ܩ#3������)��`�?�7��aG2����/��RS��'�϶b�-&�  �!��b|�Ŝ��M>��꽨�$B47)`!O�n!�K%��f�o!km|�F��:T�_?�ç3�q�Å?�S�A�o.m��RBRXr��TY���O���zU��o{�������\¹U��+u���m.쭔�P��״&�\�Q�1��9q��k�"�rN�Y`��IJ��]�U+�gB�?G���e�³��>N�(��+*���N�"�xO�E��{��9xY���g���b�����y�;ŉ��欌�z�5��hX�ѳ �ѽ��|��M��`�gqsW�)l�{�'���m��dR�.1h�c\F�cA��WB���vrY�-2�K�󎆁��w�?��N�:���c�
FdO'C���u �}�֧M+���޷{���g��I{�&���ru��۟���w�p���+�t�~����%n�eB0�5�}y���c�w�-ZS��Ί�#��r6O�tr�/��>�T�<��».3/\���$L�y��1����RtZ8ݚ'kK�B�~'�s�Jt6������}�-B��� 2�#A���S��Mk�ǑkڔI|"����'V����<�ל��fݡ�Ja�V�W��"[99�!��N/��n�ŝ����r!�������аw�a���I�c�?�}/ܝ@��oF.�����=o5	��L�j����/�7)�muYRn��g8��c)^/���<�q,��9��$B4�W"��9@s^37���K(?e7��˞?�!G�ͫDLI�m첼8�8�d����m�ƙ;S�{���k�Z�c�iAб:��ׇMU#u���wG^��}l���'� ���fe�ێf������$d�?�N!���̓��F-B�����qY!��R�v��M����b�%ي���n��|څ��{�ϖ&��^�\i���&U�l�А��R�S�������.c��k�#ͅ6�)�Ve��[�/w:/�������O�z�f����}��}wV�ïp�)�����'<���꟨ż���vk��u�N���$���E������漅/f�:k�Y�5��U��dk�z��I������O�j ~F��;V���.i��u/�s��c,5C)�v��cˎ�P�«{|��c����k9�ە�I�[��C�K� ���Ӛ�r�,��A�i`a�WK"]S	'��Fa��_1�M�! ��l��+}�v.�,�9����jx�g0By�#�T�m���AC���s����Y�k.��I��g'�	l�S��Z)[�jm��)ɻ���ۦx��}ݮ�}��v�_���2�b_��}4���C{�o�}��ɠl1Wu��2�&3k��?޴����m��[�JB�S�-�u.���>�=�{�%�UKQjI�+��z��m�3͍���$�Wկ�����;�A�Z���'-�uB�r8�;O���N%�����Q˲踦bl�؇��'�5%q��
+O,G� r��0)��@��$oy��G���3/��j̍�~�nb�o���T7�ww��?�SH#��)N%���/���m܇h�c�C�uf�,�!m���gwN��J2�ې�h�{��'��B��+0)f7~��5��^�?�h$+y�Z����3<W��c1\����9fdcT���(7��侪9/!6�G/���Q�M}��ƴ���C��V4>���D5YQ�H��*r���j�j[{�r0�2�q�m�q�3T�vۇM1��C�xA��`Rٓdx�M�|i��,��mJ�E@t
����5$:6�4H���tL�.�+X�4��$ލ�d?� �&�g��t�^J��%ԣ]6ɨ�(�}|k2{��B�pHݹC�O�]�[<����0�]:&�1ԵT��d���,��׫�%g?�/�L���ة>I��S�2"9�H\l5�11��:ȘR�tt���՞�-�	<�V�-�Lk�h}\�6����e�fm��o��g�)��°����{
��`�HL��2�$=r����Q���t�������0>� e��↋)xm�R�BDX嚜��V�+C,�MO1��Rl������;���)�e���@�#��8;]��T���Ve�P�!��/J{�B�Z�v.�7r�5'P��h&9)�[��B�{C��mOK�١_��ݗ�t�d+D��_�tz�/����D�/��K��9�"���K�Y��SE� �P���#����q�/-F�̓��T2�z9NgD�M�p�)��j�#��ź�[��ts����*���!��HZ��h�a~%$'w�c���|�E%��"`.�-�� W���Y�Lo0︽��倓�e�����G����]��rz�E�L����}=����vۊ��lu�C����m.�0�-r�����������]��GG�}Z��2��N�-Z�1"1k�m<<����߷�u��1�lIRq)>���ߒ)Դ�4rT�e�%U�ܡ|��0i�U�^�,�����&Nuˡa����૰���s������hQ2I&��]��q�����9��{��T֋*��3�8�?O�Ӳ��b�
SHw.^i�^��X��/t�o��|^� �M���ɰ
�ﲓ����-�k���X�Cn���(�o���6ȫ��ŅC���	�-�ZG!�>߉��aOF�<���Eљ�l���Φ�A���������Fڏ��C�\A&媩�L�~�"�����o���~؋qܶf���rV�Yo�aR�7�nL��@_����!h�!ي�����U¿ �EW���|G�+�m���Z>��9�J�
e����{t�����nfJ�)��^��}	i��.h����������&��#v.�F�減�w(�_�@�U�S}{mr
����~�.��C��V��:�����c��4�n20�*����!��5(g:v�ؕ8`bb�NI`����W��W�B��3\������4�KM��Ajܶo�����{$���y1�|fÞ�:��_u�-��������봾��JW�@����G����ҟ;>l`��
�"�tw�i�F�X7E\�;j8k���L�-bI��,��[E�O��HB'?H���ڽP��������&j���0ļ\$���!o�2�p�j��5/�p�ڝR%OT�H�]���P��|��g��X�8�`��'�s�1�U7vF�1�!��~�৽�BHkwlG��/�5 Զw/���\�`�A�N�AB���^����FY�-�^�ܗV0I�z��n�*�.��Gk��u� ���i�p�#Z�������GYZ}ZE�{/6J;��`�t/����|J_�]�޺�s2FB��{CBPq3#��SJ׭}�K�H�9�;
N�e��)�M�vn��ព�G��ۆ��mY������>)DՐ>���{��L^n ���dᆻ�K���+T�^~�]��l�I:�ζe�#C���
/�Zm��J߹灑�CS��6��k��`�)>��9�G}�n��xA�.r���5	Hku�	�+W���W�Z=)幛s���H 2&������d�r�&S�P���P�s2H�70�Z��Q��l����V��x��I[z(R��]�pSc�q�j�1ȃX�Ü߶����/�h�6�}�%�I\>��a�_:��R4�-���LIWј3ug	�2[��Y �N�y߉�rF/����bªt~���󲇇����"&	!s���m1����hi-��E�5�68^�p<�`Wg�#4_��e �EJ~��am��䵥L�l�(\���U)�o�m;o�)��������{rw�E!��#��W����C�q7����@E��?O��l�[!uH�ʺ�N�j'��t�1�~r���A:f�G���{��y�l���P���R����Ͽb���D�N��/��O��e|���"���x�%D�Bh����������ڱ�6�.�l��·� �,���Q�d��C����Ptp9
����\t�����]�.�ו]���>:W��n�$�nU"���Dd[g��Q�c��:���>�_mIb8��,�d[�m!��֭�����,LԬ�plK�!"i�|�p�?E�ﯢ������<:i4��V%O��>�%�Kr��/(�9��3o�B(�'���Z�ZL<]��
:��HЙ�w,;@�U���!��U�[-��N��Ļ|3O}�a�aP�؜К����m�宬��xy&����~�3�����p�\ߴ�����.��[�,u�%�4�r<Т]C��4��$�V2@3f����'dǇ��uo�Fwv����,����J�I�M7�R�R��2(�"x@B~x�xOX:�(:S�7�C�;'7��ET2�c��Br��:u�mUU�J��۴��7�	�Y!L��UGg�2���S���޷gvAz�%����b��)��,I�V]��"����43��]��%c6l�8Ǻ>T�=�W�}���J���]�[w WZ4� �L�T�@+�.�:>/W��Ǡ=:�Y�,:����|p��P�U���/�����<O*���=:v�e�t沰g�����>�	h�a�/NJJ%o�G�~�G�C���<�06���-S���*����8ʂQ�N�^Vfȍ��*���$D�O�PuE0�ι��c��Vd��=�Y�b�)�OC�'`��sp���Ơ�!F�~�| �,�V�H�7ss��9B�5Y�k����V��3���<2�j7�)�SQ�Y�P�.�w��|}�̤p��}��o���Q�(�%^�C"[i�����V��O�KJV��3���2�J��(�����Jᓆ�q�5W㴠���Z7V-6v�b�GXۥ\���M����EW���,�����,�?$��C��
�`�f4ܯ�~m�=�t%��BZ�ۜ��p��6!6�A��%'�o�g����1<ϱ�؟�{w��>��,�����[��H��Ϧ�TM;����A&��*3sB��&>og����ur}���W���	fW��XI�h���Y�n*�p�N��Tyͺ�s�=2��t�`h�j�p����Z��`�����)NwuuI����
m��t�(��}-S�����6�^/#��'��M�s�vO��X�?D���4$#�&O`�a-Y^P%J��P�����'"���־�rGtBa��"К�
&�e�g(O��)�n�1�R��4�˜��A�ԸH�$Y���VG����j/�2E��w���mE?פA\�\��=�E�U�w����w�@��o�1Q����/���#��|����=:�k;BKN�tt�C�4׮�!�"<�k�g�BX��Hh;��ޤ��ۡ/!��
���ZS���a�8x��yq�95g�s�[�Z�7�U�aX��_����"�7�f�b�5:V�s֮�t6��KC\����s'�o�yX�u��RG�$G�*��#2@zz܄��4�ѩ!�aȜ�/D|���W�ݹ�
}7ܚ�0'�,N���ݗ���YY��1, ������o.O��V/�����Ҩ[�����w�^�U��_CU�Ù^�	UQ�c�~AG6=���$��
��c���F����_z���9SN��Y�jb,.��1�O�QŇ�8)t��iֈ��g�0���i#�O_!���I�?�*���\	-�F�䜕���g�~�v)�u9n8�D>y����dQ��X��3h}B�`��0�=�sm���y�4���}�._6���w��5�u�Ɩh������VIB!炀C����\��2����=����_u���)���-��,�,^h�:����!�z4�$)z��=���@�����z��IUe��|e[d�7ن�|f��?�����ґ��`���_(!Ϳ�H�8l�;�lƿc�i�j���q�q�I�K;�>vb}����;��~Aת�z~ո�V#K�R�@��o����(���%��;�q�?)��/�MPҀ�ޙ��[��r�	GI����1���/��n�/{E�H�$�����Y��@��-�����^Y��\#�;��%�	u���='�ŠY	�%,P
g;�η�fd��D�$N�����L9T�Ԁ8OeނB�;6��Ɗ��������G��|�dk>h6��"J0i�i�-�@���qomlB ������[���RԦЉ�xY>�?z+\�������{\��g�gvJ�=h8�+���<�GO|��si�ӿl��f�q|�~i>uJMYN���w�c&�38����7� a�tl@ֹ�*;n[� �<���p��Zր�ThOc���g�\3��騭���e��_�#4�%�q���b��$�ۡ������=I�eˬ�v��-�J@��&�29[m�9�������ԑC#��;�S?��rVCN0��}��-wv�M���eY��q����V�QSf�}�������R��LY����󃚩��n3ތ�*:s�!N�Z����`w�R�WB�JיR��1�k�t��(���j%�H��r��Eg�~Ϥ�^��]�MuG�_o���T�R�2�x�ܤ��x2���CB�,�&��P�^���H̋5�"��� ���%>k'���F'�t�������|V����F�~D+ei��K����`0�Y?-'��7y����z��k��)w�eDy��3d���nkJȸ+�Ҵ����C`Q�|�#�Η���J;I������WA�x��Ń�"������Kѹ�ꘆd�P����мg��̭/�_֋�b|d�������w�~J����n�m���&/�뮷fbL�
ueR��6K�����˪���t�n�ѱg���64��V�m��'6T?GG�9<��F��Y�|�||Ӂ�bB�RW(���Ts��q�r��v�v`�\�X���۲��������f�VaH��,Ƕ�_ЅN���Y}bbZ�s��1�y�����E��:r)�I��4��Y���q>���=A���"��W>���6.5*�|�F��˄$�C��.�N^�R�{�P����G3 ��[�|M��[Ro��ODm���ͮQ���T�d���&����r�G���R��A��.)ֶ�y�ȃ�0�3��
be]���� V�+�m��_8`�ж�����_n.ה��ֲ�iSĞ��ڪ�;�!sF���3]+����m.]/g�pR��hF�;l/ޮ��@��{U*[�0��Z&�E���?�ϧ�u�a?!)�#��E��b�~�hI��j/E ��N7UP�|���%�z�&���iMM�W^� ?��Q�FBaX���ȼCY8P0�Z/�D�|�-�Zjy�5�!>�߁���Ȁ��m�R��Ϳ6��~��G�[�9�����;��T�36�������[;`G���9���yk��m��k~z4�P�9��f��S�f�k�r�I=X��L���%#�e�����~���%��E��0�����Q&E.��U�|-鿰솘Oa��n��-�����z�N����a�Ȉ��?+ �	�� �߳���~(�t�Q��H[�S��I��v�IΡ}�oT�c֕���X�o�}kb�Q���؎ǍJ9:.6�֓�:�F��<LN�R|�Y�v���Ȝ�K��=ڣ����gش��|ճY�Č�>w�Z�9#5P�P��Y���lrM���|�Wڢ����<�����N�>7^�Pi��/ <�˚��bF�p=��R��;�{eǘ�o�$��7`Y�*����ly%\�R�;�k���䬜�m��Zt�'}2����E�>C�����?υ�k(��q��*���`�9�ٞ���Q��:'��|�ϐ�g3}pt��NwX�[A�ʳˊ�����t������D���;[���5"��'����nRV�>�U9hˌ��\�sV^�J�w9�y�l֩��f��<�G}i�f�[�e�2�s�����`g�q�N�j����g[��M�m�]{S�D�B�U{��֞Q+��b����������u��>�u_眴�@PY�g���Q�>y�nc׎݉ՙ�ʺ�����ֺHR��M�,�����%����I�H���/�1;�ݔU��ٷ���7��;�@���R\v��%�Ƈ��	���*�$k��^+Y�M���H��}RDfW��jcz�a�z^��x�%�R�B��mn�6�I=�l�~	s�O���j$���_�3>�'�8�w`p4�[Gӷ���&z���{��}Gƫ��`�R�`6@Hb`�p�]��,G���]�!.���ʺ�9M�L��y����[RM�2-F��9���kʡ������M��O'���5M�M�`͉�h�Ss����@ߝ��i߼ǻ�~����a�'�۞9�6g�0�{�? �T��������[:(����o�;�T��ԮΒd���صm�(r��l&��B��̱~����A�����ln.�������[H�����Eݓ�5�GI���&`����g�A��R�|��>�K5i8���
D5�,_�|�YԊ!�4	m���ӦTh�<VAiq`1zi��^\�����)��5�{�NY�ql�$c�M���?r8�N#|閖$���A����*��oA�IԏyX���\U5�=wg��|5�;��L�M�#�+3��1�U[��}z���n�\]���|��⮩+㷟#��r���|s�ɋ�tM�-�_N��u��X��1ꮚ�$�b<P�	� m"A��m2|������g�'��E��K▁���%i�E ���w�Q;	!��&���Y�L0�Y���Y�v����`����GGdz��Yg*�3�x]���y	j�zn�t��2@�i��b.j�>ݫ��t`�[�L�ӽ�m3�Q�csj�J*��7�&���ksˌ|�j��돝�X��,n�K�=tDH�UҔQ:���/#��>�(DL�t>�����7>�O�]^g
F��k�
:�����k艝q6�wD ����*[��J������������ƫvHΙ�cV1(����̖�V1�_�`C���Ni܏��P�nzO곐�&g+��J3县�B��d�w�>�z�ylu�:�R�"�S2�/6{���yw�^'���]�E��9�c���⧝��&�n9K����z`�Y�B��g���%����"K�Q[��Ŭ���m�UM^����AD'+�4@����V���w�V�J��?]�;
��4\TV*]���3xjnxGG���G��+���S�����nТ��Ҧ�$�BI�G�TV�`]ct��B6$�]��A}n���<*e��}���$0��@�A���X�§?�*Ҥ���Gx�vE-#�������kk�	g��`�o�� Clً'�-2'�[�4��&�URQ
u��eH#U��f^��[,K��5�/�VԜ]�2V:���#�{�[���~B� /\	���� !�5��ȣ�������;��7�m��d��9o�ID�?��:�#�W(��U^�f`0�|Z�L�q���ku�j�4UJ�Ӝ��-s�{%f|����zmt��GM�0Tu�_�0�
o�'�'��df�X�'�U�>ha榬��a�d��!1�RT�k��]�144�w��.���K�x���,\t��߷�6�?�.P��H��}�[ �f_7���?Us�_g��k�ܑ\��S��('T��ѿ�[�0o(�'5�w�܊'��	j��U��|#�?J����spey���Af����әؐ���?�̝�-���+�;a}|������>P���䏻�gߩ�$V�>���%���Ǧl/�c-H	�>5j6�!�#�V�es�'w��jM���:��\��4l5(��g,#��0��B��{W�Q�	�j����\*�>
j�j�� F^H�n-^G�9n]��?0�+�������õ���+�u���
9)�b�>0V�jŕ{�,Vƃ�1�T��2}/�C\ZX�v>s2�w��0���O'�ՋId��)�ؽ���;*hV+L�=+y�ɲ�{w�zСgM�l�g��/�\_[�(�x|��Y2Tu� �5H'x]��NC� 8vx� =�\��T��?&�2ۿ�vT�
ղ���ZW��Y�qC(ȫ���~��+ �|'������h��EX��HԀ���Ԑܻ��o��aL����ߴ���]
��@���(lW<ƇO׈$�erƭ����c�"{G?m7�g;��Lj��3����9A'��Ś��^��_�������r������e�#I��)S���RN�4�`"f��Dn�6�m�#p���|1Ԅ
l�­���lVj?|��"���8��4�p�6?����}r/������D���8��@=��2w�:���w|����A��6ϲ]�&�Ⱦ"si]H���p�VzrϷ�N�C���+���l�jC�[DK��*S��D�؜�5g�暼,S�eZ$����{�Bܤ\7���A�����Ъ�� Di��r������2Y~��L}�����n�� UN79^�k��#��mQ	B�OS<�Bz���� U{,cܪ
��J��U���܂�}�[�2G)����1"9�x,�xL%9�<B�4(��^���"�]�}M��S���9^��܀Ԅ�SLڵpAX:�=��'V����
��=ˮ��ʏ
�A'B�q��,��Ke�#�j
s�t�#�L�vٕ$�`^��@����,�k��<'f�L7l���Sή��H�CW�8�q����ܚ4���>���N�v+�d�6�R2��Էʶ�fj�Q�YhV0ŋ���iVǛ0h���t�\���3Q�P�_T�I���*c�ם�L%O}F�G�&�e�zwJ
F�M����q�6~o�{2��;�J�SӞ�.���ݚץ!���?�����*Wf�5��DE߉ų��S�;�{N/l���F�y�[��>�p��ț�<m��NL���饷���Jdnd��`P-�W�!�}�o� ��x=-�̋����^S�=��W��>�������*l2y2�}d�9Z����^}�{�H	e�/�R�����w�?��dVJ�B�k�����\�ߣ��'Rgr���v2�g�����	(�ag\GݞϻF���$ɐ��F�؀�d����b�}����L�~��I1a}ޮ9P`币?��]v����Lr,,�D�#LO�Ԣ����B"��i`�t宮S��	��
e�B��
M�ܷ�z��!T��������;+��KkV{ƿ\J�o��v{?#D 8�����ü\��\� � 4���wcŇ�,,�t�+,u��j�BOҰڏS�������<�K�yF�"�A�������W
h��\9��#�9�����ٽ&�(�+NX�C�V��bfv����E���3�{i���D�rƀ�e��D�{�ltv_�:qJv�C�w�����g>�{M��C������H~��ZM`9���Ws#����|E�ڞ�ZI��F�2CGD���_��.��v�uAJZ�")���
x�%�z�1ԗCwW{)��������n���@���?L�Z�ea�.Ł���%�j��<�+k�����w��*�?/���ll�����(���gBh죺�sU&{�yo��"<�<�+��+�}ú���I@�f;���Hk�����{��`nB<�fl���u�EceѺ wL;��2��hQ0�;y��<�7��k#y����ϗ�6�9�x�ӭv���x�6Cs���a�G�r���z���JL��Z��x;;}�E<�r�c�7���$�C��%e��R�H]��YҸ�^|�v��H�iVq�5����Y�]�r��4�ߤa��s��ˌ���+��bns?]�뵣׉��Ɔ����g6f@��P�M��ά��}.!��ޒv_I�wy���J�gr��TH�
tT+�S�w�͛�zݿ�O�����N�\ԓ��5Rq���J�UÙ����Sb`l�E`�S�ĩǸ�PEFi"b�pF�GD*¶��\P�MA-�U�T��N�^�Hkt��[��ߞ�-�����GH��+:,����V������h�r3}�>Z�������㫾�Ǫ�Lg'��w�G�5Y�*���q5�;z淾vx.�O���ĞQ�#!$_��dq��{P��P�Z��ʪd�B��ې����rm2J�mvE���t�����&��@��	'0�M�p�(; ���n`�g�� �b��y�Ku�����<�8|\��ʼ_���������mQX6*�k�AW����״é8�exǻ�*Ҭ�SW�7���#�e<'S��갈���r�ǜ����ϋ�
�Z�N{���׍�Ӊ&,'|�����QlKi{"�����{�7��w^օ⃣!ɪ.�}AX���	�s���eR�p�z�~"�l����4�u�|-�i��}ee�����pr�^��n-���ڤWV�п�r��A��_�Zo�k�`n�.��p:�Xo��.Xޤ��,7�st�a�~�X]�"�@�#�*8{��6m俣�!:ǟz����
]��ɖ��j��ɿi�bL�O�����By��eV`�z���g�z=/^��T=�M�cIt��4毓���jޏ�f���TD~���ʤ��>���� 3+��2����/j����\�qF�����!��9� �A��),�]�Ż)��ti�n ^N��y:~�s6��lWSA8������m�/QN�6*�B�osS���š��;߼��p���ʨ��`b-2��c���oy�$��j��si�����e���'1jLKa�]H�3�Ш���l��;��3���\��\�cP��_���y@c�0�S����=����v��kӓ:�Է)g�쳙����H�G��(���?Uy���+�����hCՋ��������I�҇��ϔ��ʕ�1ۑ�P�vX�"�64T^���I�oy�@�a��m�cc��N�?+�g��J�9�a�p�.WP/k �s�#��X�!�<����5kG�~}��]�T����)�SF��l|����FY�l�����4ֿ0��@=�@��5���n V�炚���G��	N.�\5�N���h+�G�q4/�f�������@�M�t�唙u�����!�=Ó^��������)��l���#�h����u	A\ɛ�k	q�r(��b�q&ٺ�)�5��z�<�ҩ����e?�2����
�7�Nu).W�1	y3�T��bM�IZ�0�n�'�K�4�C�� ƞq�֝��({��h�`UF_�L4;7�H�f�e���Z%���[�����s�x�������e���9\}���/�.g0�q�Öxo��ڬ۳�����d2��[�.� �]��M�1y��a��9d
-?~����Pa�'�YI������f�K�~3�St��T�O;Z������:�Κ~�� �������A1�ק_gg��Z}���j�nW���x���p�/w�^�8Q9�ǳ�}� �_��a�-"hX��湣!���E>�3_?淵��G��&2D�:��Jr���R,�;����V�D=� � b�U.�6*�"8�?P���0��YQ�\@�j����zWV��f�:8�5�d<�Ӷ����}F�	>�&%�/�zH��"�G(OE�JEސܣAhLהz��	�$�q������xi=3����/��in�.r���}�\S���|<�G�����Y��Q�U/��Oml<�q����>p�ԓ��l�4�|P�EfE��=�-�u ���E�)��ʯx�ߧj��1x��j��2R�$哦��"���^x&��5�i\�-��<#��y�)��	�����K����!����RXc96g/"M���K���iWt���y�W��z	�ȕ� r#�W��*�|�<jh&�v��d�r$���)�'HHLb_f�����P�)�&�
M|Nl��w�@/��gg�P�[�l�Bm϶M(�I���R���
�=������eS����	��+���kb�A]�͑rHu�c-�
L�nb�vu��>FnD��]C[g�HW�m/����������q�3`ZHM���Q��D�7D��w{oS�H:\{��e�-��?�~�vt������i�,h�q*��v��(l,��ޣ���`���Lo�5�OB��ˬZБ7xO(kP��ָ�^<�KB����);4&˥�kkr����r�K8����5=�c5	η�Yb��hk=����
��Czf�irw���m�E��1�
��Uh����ɻM5٥�ȟWe���I��0�<#|)zN��ERԊS's�^�}n�����I�J��50j�U�n�����[۷Q)�}<�Q[�V�؇�hi=	�UH�k�r�]^�R0�!���rNAY�;�X�嵉�. ��Ne�BҠ�Q�ӋH��s-]½�N�9��"62v�V�g���6`��s�ۛ�e��dF+]�DŸ(ג$"~�Y&�du\�>�-O��\*���W��؂�#*�Y(��s�.��rb�2D���[2�w<9R���e��j؎��L`�c�O���q��o���A'Ǖ�0R�::��[~����¡���=�%�)opnً)K�9�[r�"
�_�S�P3���S����j(Z��ɔ:d'Q���F3UW^~zY�2ȼ����+%���"ʩ1H�ߖ�ƃ�ԇ��
���*A|�\���2o�mm�vʵ������JV�gh��(o�~nڂا��[��z�����5��qד��ά����2p��nӻG�������f��t9����ک���ٓ�Bָ83���m0�U��!zDѪ�������-��v�\Q�G��~����m�&�o\I{g%&GԢ�/�FMz 3sn~��?}��%*6
E�U���r�킡��25|�~����;�?��'���?W?,��$X�J�q�4?��r�v�j����i����{��5�d����@�Q(qE1s�Y�|ƴ��4u�כQ��)�ż6��Rsi�3�U/�c�%?�/�%(�,��}�)}縒b��۹ݓ2]hztPo��g�����]C�g�p�,�45�k(ȓ�i>3"�l~*�[˿k�v�{c�ݭ稺�Db<��eK�C 5Ԣ-���T�%��׹�BD���J�`Y�3���R$������#�����sAsu�[����w��2�:�?� ��I��5<X��h�:�/�O4���|H���!uKq�l��p>�:Z9�6��T�d���ˬ�� 2�c\��1�}@��[߁6�e|��&;��wX�������2"�eu�K���s���#�2"ף��R��@
i�/7t� Z?'Q|�*��g�e��Nwz�,I|)]JZ�*!MW�h8�ѯK[t��+�b�&�j{�`��hg��!]ʰ3��9�������p��9�̝�����%r�2����j�F���'
��,3SSi_�TЯ�%
�7��iy�������~�3��t�]�;�G�YZ�bs�����7�-ML`�m)[
ݖ�:��D�v� . AEմD� x,M�Q�����r�3}�$E�+��4�VG���\]�r<�ۓ����°��GUJ�����Y&>�1dm5x�	D�c��*�b�K�o5�> j\.Zj�CY4~�`�u��Lз%vE��au�t!֣�v��˅��LJv�3����8U�l2�q^P�(o�L�l�/RqY�ǅ���Z��,�+�d��{d#D>#��
�X#�P*�<6����bw�ֶ1��-'���)Ig���DI��:'	�^�Ň3�Ą@��	fe3�i(�N�m�qU�ѕ�z�FW�+x\�RҌ�l5l
�rp7��� �v��i�8���:q���ݒ��f���#ٺ��d��^�]+c����eK�3ؗ�(�Ӫ�/�/Dl�kteOp�4����Sl/�R���5��Dt]^�Z�3��9���ښ������y������nD�("Ϫ�h{S�<u�qJ$au�g������Q��՗mi��9X� �e9Yl���>��R14n�~�fo�^�\o�'c(����JԦK�95O�B�a��I��j
,�ࡿ�9�6>��M�ԆY{ Jg����~���X8���ؐ�	�:������ЕT���m:0�uPKs������7��*$�
H����t��oE��9ƍ#���Y̸?���4\�#欒=��!bDU/ �|\C�:��(c��s�-o���pt(��wm�͚N��]o�XNN�"yQ����R1w��L��ݮ|XԻ����#�����b�����탂Z<2+�]��8��aH["f�|L���!,�^�2->93����~S����Ņ0?���J&�ڡ�A� ��p�c�=������݁P�_VXL��4��ni�BY���0�������L��PSE6�w l��B�An_ۊR?�+����:�`�����o�Q��V���}��Ѽ=?oK�]�:l
���T�H�������Ǖ(+T��;r|�����wr1��_�	�m�^	)K��-��$d�^�sϋ^�@kgo])&+����"{G�	��K*�xy����A{�~�x�_��a����niiA����ɆQga+f9PfU��j���L������ͦlwQ)��^�\���Q����&k��u�1M�f��������}b;�ըm�&ήiΟn�k(��*��ߐm�i��bH�S�G�H�x:�jS7������Ok1q�t?QZ��U�Q"��ꐺM�yq�R.:B5A������[��c"�����,_Jf� �r0c�r�`�㧡�� ��d��a��"�i�т����ۻq�gK�c`oG���ة���Ϋ�^1�&&�}��!�`����+%
��9���K�$3����I��s����6o�I��lW�:�3��{�ͪ��w)�n�/�Yą��l���WϾI�y��Qޓi.u@�D-J�R�9#D5Kƕ����j��2��muy�}�Ov��\�u��u>�|�y�=7�ov����;�m!f�6�W,6�V�z����U��z�����o�ge~X��b�2$��O���p�OS����:��?�[۷�KΝ_^�!AC�y���p�WX \<x�������t�NcNsm�&�ȉ*mҠ���"2o�I+�������a����	Ue�ץ�8���{-v�MG��ʘ]�f aeRݺ���f�;X�	�U?
.H�\a���x1�1���;�d l#������3�\��D�~���5aǆK��i��%v�q�}#$to0��w@��K���G����{G�2#�;<[ў�sI��'�&�=J$L���FxL�OJ�;�vWD��^2�*6I�C�RI��K��w�{�.�_]�{gB������4�+��b7����S��V��o�Nľ�/`�q*�g��#d�=5�7�l�+~�H�T������A�����z��.j8-0[nJΑ�)�5ә�v E�?e����=n��4h�Kk�'�������@��^�#eB",��eU$x
m�L�h��[<>��g�f4��HK��V��Ft�Sw��๾���ݞ�=N��G<]3�����0�7�q���.#<����6j�!�04a�	��Ex�V�"aM7��gH��J�H�(��w.��Qp������ 2�lz���������l��n��� R���ף��/+��&��X���*r�6���*�L�g��.�f^2qn��+���0�CŽ~߳ν �'x�����.���EU����l�w���p�o;�/W|�q۟����S��D�Rg�(�$�}�e[�G��סM����Wے܄��b�H��´���ڇ��zSD:�@��,?*����=l˚�+v�M�S��<����p<�W��1��	/O��jѸ-XrkFN�����aȕ\�_Ӑ�u�6W��ji(��ٲ\w������(�4b	N�Oo���N����i��j�����W^�����!;BČ�qk�;�R�c�%>9���n���;{W��d�U�����޲�yzmm����8� "ֻ�~F�P��x"�D�g�K��6�n5V)>�T��wJv�����CY�H~��O�N����������h�)c?;��S�� �F��^O
(z�}�o��K�&���塻�mќ��uXͿX��\�K%������@8h;��a3t=߽*wXMK�MW�7�8�I%�̺> �!-}�3{�m��A/�8q>y��fP��{Q���MKX���Xb%n ��@��$�.��tsA	³���*��`U5�&�C�/���5*�v��f��%TTbJ��c[ƬyA��6'����X�4��yq�.�<m��}X�k��%�ދ��X��oP����{U������uDfv=�C�k�)	�Q�g�4T��o¿G����7`�t:[6���˜��!Սn���2��á������6�)�㟮c������6�89& �N���	BV�I�(����nI��;��Ӹ���Y5�ףWw,CY�:��yqۙ*tX$_���Y��݂�`q���~=f��R�O�@+),��U�h�-kW���H�;/��^D2��o_M��T��U�:�A���MS���\�����ڰ^��10�����Mj*zr��������i�]B���|�"ˬè<;�f�k�E�P�ZciR���d����PI 8@��Ր�:1r;`������"�����f�ϼ_��r"߷|�H�.M.]x��8�?�w���rP��2��<�J5�������ڶ-�f�e��������uO���\�s� �,�	�y������a��l�6b,r7��Bg��	��l�乥6N2"�&!�VB�osM�`�o<�3A[l���~)��a�E�c�H���=䲷3oI�؊sN�9y�xd�[5}�o�	�r�&����g�cA�^tn��� Sݫ�����<�֐��8����m+��������Fп�a�?]5u�{(��G�H"x�ݘ�T�/�6_�}-&I��,���wߔ�i~Gv݄B�ż��� h'ӓݻKM�^�ܯl�h{�9����6�]o��9l�����
�<'��5.����O?�)o�G��u�.�"��z�)
��e�����0�+��>7)D�5x�g�/�-,���is�����=1TM��ט u|�;i�I�^�&iz�>j���<O*`�RzXJ��|ӎ���x�lOif�e}Sa��0�(�H���-"?@s�.\�,�w�yf]��@�V>�O��2�8�j5�f�pxXȳ&�Wm�Z:�� �	�,�C�/�����d<���BO���i=z@�.���n;���1�@Ng�����F������������Dl/{rX�^�e���������Hul*�y����1��N,`z�Ļ˓_�&��tQ6���O2�ޝY�}C�ɭb��+�f��}OUjUu�gyC�ӯ3ռJC���o]�E��Ꮧ�1�d#�fބ��p��n�ѯ{ Q�7٠k;���ܟvJ]�B���9��b�7��1n���`k�|����&�<>3j���&�L��(\-.Gp��󖎒�P\,��Z(�#�1�x�TB3Pf8($*e�x�ʕ#A�v�yy����hmNY�UF�m�,O���ɮG���e	��f���X�Nn�r�R9��o�lm6�.Bc�w��6Z���#9��S{T�%syo>�(p��-��(�N$����i?Yں���nA�`���������s�l�{�˖Se�)�f~���0�Е�J;s_���}_��&�5��(p��g��k���<�Z�g��=1�|�o����@���ن�:�Di�1���N���P-�e�&�"�*Q�nxqs�I
�a��e}Z-��b������_��{ȡ"˹o�]xӦ%���)$/�'Lq�3UHT�l�i-���a���ug���?l#�W�=��M�}��J���u�SZ�ɿ�$�|�T��~ªϞM�1h��n����m����䣖�'{(��.):�mdG�]*�K�P֦k�=\W1)�BM��%
:��!�U�]&���C~�7�+6ڃ�t�%q��q��S}����-����]m>)d�8W�{��Xv@���^��1���<�X�OF�����KU��Sl�4h$��A��g�DKe0)�PC%T�Q˖u�[�J�}��d�	��e�:'�Rw�ӏ�Y�ԅS��0��Ɇ�7���\��d&t�P� |z	$��F �7-�c�JktEo��-iǸ��5�!8@E�R������P2��<ogE�������Ok-�7�p�&��5��'��^S�ȋ|_�*HF�I�����$��0�\����NB�����+��wP������`_=�!L�n�Q.�O�&kޭb[5�����>�~T���M|yP_���R� �#cD�D*xJT�%7�v����oM�p���b�So��:��7kך����=��;7" z�k^my�g��RÉ�	D���i�PS'O�w2z����.d���,$U^�5H��/v��4��Ku�[GH�/6P��0����EޙKi���@���U�-#�O��lV��P��!"���7Bsi�XT7z4�"m�fz��;��n��q��7�u��j�Sõ�*T"ptd�o�-�����xf�L�{r?��������Y��L�[eu��=�:G ��9�Ό�jn@��N�#���H�����>k�V�/c��m������ 3�����l�BadUձBri�%��۴х���zNҨq�u�)h�KN�?�j��^�搆Ƴ�s�1�0����>��
0Q�Ij�`�YtHe�]�� f!����Bc��������������ċ&��z�0�����q�A�)��G�ȘD� ����aE��gx��� ��#��B>0��*����S���n�ͦ��:���R�+�S2�.�\���%̈�Sޟ9ծHwę�Z���`��ڄ*eB@�W���"!vh�E����^�{5�>�.K⣥�Qzz�fj(�ट��]�1�y1�?����&�֎ȥ���0x�,E���E�Ӑ!�M�d�[��7��2w7!i�!9�jщ44p	T<�t��ɢ���2w�c{X���&{���d�6J��E2�wq���/nל����ZI���P�K��O�	%G��=%��LY�h�@?{����Wf�kzJ�q���M��~����t�+�V:��V���+6sk/�4�V�l]�=^K�Ϻ�ם�������&�����L8;fX�B��(:&���=3Y�w�s�y(�99��;y�S�bP=���M*�v6�Ku�:�h:�9x�0d�;oZ�t�����l���:"r���?�o9i.����$�A����D��H���xUO7i)*�T�V\��ߨ��[C�)ֳ4����k�_z7��L�M�.�*D�"d��بs�	����ҍ�C5k�p�Q�ѭ��[�65��@�3�¼~Dn��KONn7����\i�x?Y6�Җr�B����u�!��(ͬx�	�5*c�f9kL%uǟU�ӻ���Ȥ�X@[u�K{h��[��7��P6\��`0��Iw�u�c��R�e�&-�P�ܙ�J���#�����^�;��{ٟ=�2�yL�B�'�^e."�s���C̰&Z�tԨ�i�̀�`yص���]�Z,$����1���~����l�,��o�z4.����˺u����6�����Mg�Az��n�����$��L]%�g�W��	Lz �֬&�f��`l�}�9��ny�M�z��k��(���+�qͱ�v��:f�ؖ��v�Q3��&���;n }�}��#�m���K6o� �iY���})k�\���DdT�R)�g)�G�>�Pt���d��oR�V!�����۔Vf�����z���w(�G��h&��\�$��_��`|؀�t�^˻ /z�֚�d�6ε��7�^N/���ϟ���)\���7����p^c�.���}<���%
:6aG���8/�a�Z����)Zz�eH����Ҽ�D�˺�,%�N��8����o���F��g,����H),.�XtY-��}���2=�����*1;{A����������
��ub	T��|�0�=fp��0��[#n���ゴ��9�wvX��#͈E(a�ٗ�-�ñz��%������]u��K7���T�c0�#�M��M=֫�α�Hv�v}�`�y4pd|A��J��W
�z}�1�ִ��f@��)e����E�'\x�`����f�-d��?�Z�.o�ӾqJ�����[�b��h B�>��.�so � qm}�����wWD\���nB���5}��."Vq����=��ّ�����'.���z͢�4��r�w_���)��S2[��3i���(�6[<]�)��ޟIiHa�ךd5ƚX�<j�
jM�c��g�}+�������P��@T@1���ϳ�K\�������?G�S���K��ˋ��f�ĸ��
���hyB������f5Y�,���)V��$voS�<	p>����7`�/#=.���G3T��.vѼ^�{x�������L�[o<3���,rK����-9{�R�/��%[s���&�M����R1����9��g��m*}k"�J!\�'<��slq�Mr�7A�T��||c!W���D�f�uInU����[���7�����f��Q�S6��>ey�t�a��HX�zLCz>��PX�`bh� Y�AиA�M��~>O�ڸ m�!n���jQJ��'챨�l�޸���P����N�`M� R�m7R����H�	���K���;���-Uh�YSu����=��kE[�X���E��p�`v^�>Rp��`�~�n�-7lw��3��n����
�/o&9��I=�m����XW�u���[\%��{���;��Y ��t��������j�)Cqt
��8��=�PI�i�bf:#5�*�j��M�3p�{�Suү�^#\$C�tt���`i�B�
eNx:'���~vc��226��	c�
{%S����B��� ����gR*�;W��Ck}VP0�~�Q���#SZ���%se��S��ѭ�	��y��.'�`��j_?��P-v��Z�+��*+�q`eT�:؝۳k�[����ɤ4G�K���o�o���R�t�2��U��+_x��1pa�v�5Hc;�տ�yP��7D���f���yT���ov:|�|�݄����hpW���[�lz�!.�4b��ks��R��0ם�Vaʕ3����db��ë*$l�$o'RC��xg���4pN���&��8sk&̎�~��ö����S�V)xZ|j��ZK�g�z��9���
�[9=w�e# �@j^;�Ҧ��y��n��*��(x��f������w��R�(��e���qx�і�9�u��H��5=86-/���F�V��Z�c�G�Xt^R��!1��+Cp�ir	��5]B.�dwL�5Q����O��3X���n�Y-j�q:K��|�z����	��{��̗�I���N��L�Q�?���xbV��֩��bm��:��S��~o4���.� �2\�;Cʆ�&v��?!v�g�d��W֍v)M�^^�LxWT��KW��.xM�0�������)�'��힫���/�0�|�>0ƥ7��]-ی�V��N��<"�6�����,6kʯ��~�}��63O��� �"Ti�:��>�T�㷓G�/���Ս5��Jf4��^w`@ ��WZ\��l���`��y��U`՟�F�A� �Z�ӜD1�����?	��Ǯ�Ԋ-:�+�ᢄ�/($k�}��LY��}�i7i8��1���+-���S�k8>h)9N�-7�K�"C�XWEc�Q�i�b㺵�E�?O.�Q����S�����*���fΧh��犔���]�(�:������m+(|g�&�DHG�1����M���!,�]OE�r��F�l"[����Q� 5:Oۯ�����ά��X�w�7��F�<��!�/6��ւP�Dd��5���� #
+��M����0%��GJ��Y3��ۏXqZ�w�/�̗��f�U����n����jd���ާ��q����`� ������ƕ}{Xa;Q�@}���w�kq��Qc��g<���R�%H�)E��q�k�Q2������u!
&��l��<�Ll6p���6�(^���BǛ�b°����J�t��J���� ���#�;��P���j��E��n)�)joګ�Z�7�El���Z����ڛ��l��++�� Fl5~��/|~���<�{�y�s�CW����]M�{H���vKH�z�������Q#�ݎ�C��lK�w���+�H�4;~���'�s��w��t|o���H[+�Yt���VH�}\��47ɦ��aN�o���g7]����0���,�[]�x�x�hE �xA��N�C�2q�q~b�~�:�pʠ�ل��Z�AX96OOhhb�Ֆ�׸I&��t-^#����05� n����u%kɂ���)�D���G�
:5Էa6���g���T����<Jd��ݕh�$Q]p�ߟZ���qA���@o*%�U�/���-MR�o.��3�b���w��ı���^7���eoq��;]�}&&�ZT�M����X��Ԕ$@V�����
��ҝW�vt�	(�9``�97}~�g_���%�.�� 9��X��֘�_?�z�(��vG�+TC�n�{V'���Rs8��L)3
�,5-9����na�Y����]����U(\��<����vL��o*��BC�s�9�1����yjs����I�5����$>�"33qHf�	���� �~�1��0��f��K_�Y�V3��ߙ6�?��s��ąx���:�
���m�=��\LgwEw���J;�I�ޫ����J�IoW�G9���K��<��4��yk�7߰t�.;��W�}�gΆwc���c�DPA���i�,^�n>�U*�Ǩ�&FyΕ��2p�T���zS�"월)_t0�,���������G��R$��= ��ԯ��p1p����`�^fK�qß[��M!��1��I�X5�� �SK�-�=9�x��������H?���ϲ��3�L�m'jF_u�n���K��+�X�'
zz2���W8�2����;t�e�n�����lt����L�Un���^�Ҍ0��ē8�k�4'��v�VDFQC�O���w����A�)R�Q?Ă�������J�Nm����
���4b�_=�(���1�� �GG+ҳ�m}��?�zzˊ�4����Ն�8�)^��ۤk�O�C��7�^��������ψz�b�ft�!Y�h����4�����c�d�"��1�cx<�����+D�����3N���77�ɽȑ���V/"d�3�W�nt�>͛�jR2S������y�肬��������.t |��C$�R�h���8�����z-�������3v�L^x��g��@૨N���;GE.�= �CgW�ݰ�~f�ɧA�.r�S��Bɖ#����-�X�Г��;����m��9�h��cI�����'��;'��<�V\J�D�)����.�;��v(�a�Wǂ�[:rƈ��W��g��n������JK|��Z�X޾<��VA�4Q��O:��4�e��I�K�L�y\���QRTD�:�Uo'�Q��l(��8�椆�{9��_$�'aC����eO2�M�*���t�<zV$9����R���:�v���Ḯ����oSis��M??:\za�������Yw� �%��l���Ǉ�e�q�@|�c�G�xo"84��OgSmq)v�� 6!��c��A��MFA�]r�[�yA&G;-�����bF��f�M�����$"F�������N�=�!��X6��|��qr��eF�B�7�n~\h�z���+hCud�|"�MqtP��c's�R�u�v���f�>n��J�i�CZ��R�Z����O��ټ�p����xx���r�S�.��r��%Т2-��@j�u���Gp����35�.V�SoN`�1Q�_DK�!P�[��$$U����Q�CƄ���Yh�n.I`<͡NQ��wSmF��<����v�Hn#:��UX&�YB���<+��M��X�?�Կ�]���U��Y6��S#|�TdIV郖o�u}ޭU���羢ll)2̆&�Qݓ���ꑍ�V�����������I>�����Z�~��T���� &#��psH%sM�D�{˓��������!�ʒTXh�5.�]�K���+U�|�籍Q�0 ���c���'�%Y����J{'��C�G���w��Qwn�[�?Qa
��8�H��͕�i� ���`݆��z��E��AT��4j��B�E�O���]���U�[��GEq��=\��Wx�ǃ�$�)�@K8������g��x�uV�;���/�q3q�u�����h���H!����e�����'ηB��9�����3G)t���s}�%��w�J�*ʓ;r����	�9V�n؅"|ѵ���������܄!n����=c�JkK#�� �%����.�5@9̱�<hw��i�ϱ��z��)�-1 �<s,�\3i5�O������>�����>|@�ϗ̨�p@9��@U	�p��y��� 4����~���0�#���e�1�2~�j�5gz+Q(��{��%KwM��:&��M1詫�c�%�.@���H q>E�';$4>�]��s�(?V���
"�B<8�(���NPs:m4O<�@=���?�ml����^�6x�*��a�7�2�aq���6ϟ.�K��%dA S%fu�+N�h8��T��8�x�)��!�GpG\4=��t=ӭ{����0�с�����(>��2�p���<+O�Fq7._2*����FQ�4��qj�x��+k��Oh�/�T����`lF�A�v�i��O	��"�1�)�b�r[c%ň�fS�ʥџ�3kO@<}� �b�C��2�JM|�Y�a��v���mV�I��T��$��@E�_�=�t<�n30ʹ.�K��ޞ����=�:���X)������S��x���������?c/�hjH�F���(�|#OIE,���w��`�GhU�Qa�Pp��%���hm�r���b��UQ� 5�X�k��=_s�&`Nx��s��'��N�l$f��)�ͷ�]B��G��{�.�@ߊA���B�g�C�q���K��&r�ˁ�[j�VE�I4V�L��&���Jsr�^���������I���l�QoJ�Ks����|x�o	�\�u`I��/�ގ4�S�xaN��y�H�ѲG�X�і�xZ����Y�M��E�1��
���/�Φn7�8��{tt�je3D�&�7�k0��~��"H>��F�f�\x���"����I�˟�yӽ1�"|�x����|C3u�J�QJ�R���h}��BN��ptq7$N��g??5�i�O���y��T��Ǭ�]�~Vx��n�;jV�c��گ���jH+>(l���{QO����y����7h$�a��o=�|m>����t^��E̙^�-2�_��n-� tum �(8���G�<�Q+I�c�s��F1���>���$
±~l*�$n��l�c�cw�}sڮ���|�v�~�)B�)���iY��QeI6~���r?֐����}���믢���3�.����'LJF$9G�LPl6*�k��i���ׄ�Zg�Pd)����]���V��$5r�����V�t�{{C!����.<���ڪ�L�TæD�-��~�6�P��e��e¼#E;�-�ǭ�FV��#���c��#��x(�Ë͜�����$�����L�{GBD[v�VE�߽8�Ғ<����s��KQ��P�#��t6�C�^�6��ф�;�t���|s���Kw:`��8���m~�p���04���;P���ҕ7��O�o�e�D2���R��L�Խ)��6���8d�u��g��b^��b���o�PY�5�+�+5��;�0�)��B"jzV�n�J/�9�
�x��HY�\���V�����1g�_��ZmV/}L�CB�+���N�61�6v!��V�^ڬ�|�G��	\��2�l�'Z�<�u#��	M��ڥS��d������iJ���ֽ6&��^F��+�2�ԕa�k��[!�՚:D�A�:����m�H���'�V��Ҝ)����>�@Yw��F�
���Z�$겺��7?y�j'�r ����Y�RI[��p�uA�\�r-[�`�ՃE�g_pd0�4-��Q��&,��B�C7�ƒ���2XJr�@jh��W329 s0����f���O}:']�õ���'�ʋ>D�$X).��N]��@�ܿ�;c��Tn�F�J}W�F[�[&(��B�$O."R��ܴ!G��{�+<�\P՟j��E�_cI�U�ŮP��*�@�C�Ư�~�4;�ur��M�Qt�~8`���_*hm�~
���;��z�gW~��<d����r�ު�+V�z�~{��$���U���u�M��Mު4��
N������x�XZ�W1X��Lޟ8'?TG%���E�l5�ݸKZ�X)lߙD�d��=��uh�9i�Z��<�|Ն3��bUs��U?̞��|�~��6�Ⱦb�7	3�o��f�KḼ�Kͺ�;��.̰^|��SW����|��4�����ƞP+�ʉ�*�*s���/�LF�˨ڌ5�h`�Vɘ�R�C ���*�Y/h9������z���O5U�m��0�yx�.�M״I��b� q�:���e�<�g����,��e~��X�Zp��i�O��z�]�V�Q꿣J�Y1^���m�ߥ֗���2�5}��J9�bf���f��R��I�
#ujbr���t��w!ƙ$�<�4��G��"EC�dJ�LW3 q��h7��3Ҁ�$6��J�9f}�<vf\��6�Hw?e]Oa�����]�va�f�����m�:T�$M�½;���m�v޵��N�Ɣ1�>�t�m�������}L
��O}F�PGyDm������ �)Y֦!��C�7�-�̋�?�<��8�R�O�dU��鯙������Xs�֬�y5ñ�{���������a66Ϳ�_<��Y�½����]M�X�/��{����§�Sr��u����� Ӈ|6L�y�,>���m��x$����ahF��w���}�`�Ж�>(����G�C.���7�{�ZDY�qh?������m_j@�O���b4 r�Ơ��q =Pf�5Y���5!~ϩ��`�L���yn	��ثd%'�飨Q�Z��+?�YA��擐%��h+�(�L#�N��a�݁�)�ފKm�~?t�w�d	r���z�=� k���.�T�N����x���Y���;�d�ov�x��ݪj�1iX�Zi}D���US"�/�-6/�e/L�����βI��h�w5A8���:�C1/�s��+��:��az끮�+{J�����J���@e��������7�F�A���[��{���i�����;X��t�y��K��;��_5���;��rP{�r�
�S����uqL��ea3������<ԙΜ;u�d� ��1gӿ��&����O��;�e���&�ȴ�b:KC���{��6���3�2y~;����q\�0w�]K����mb��17�b�D�����9}5Y�p�8ҵ��bѵ��j��=1��j4zc"$i�M}�WRˑvbiyv.A.n{�)��)��<OqZ����M=S�M:ֵ�j��l�W������<�;�����"�u�����7 �%��r����I������T���4��t�c9]�^[VYSWA���Z�CF(��"�Tk�@���IM���K�"'\�ي�zffU^��y%XP�c����C,�P��g#{��%KY����b-��6>'�if�=�I�����3d8,��[�%^�wOkk;|�jJA�
?�{0���9I�!��պ� ���lr���ˆ{F�|"� y�5����i�+�Y6��:ڞJtGK��BPx��zF���C;�f�wa&�0͜z��J��Sʨ�F���|���s��RD�|vI~ۍ��+EU��fjR�\��$�_G�Ph�W���{h5���-Z��'я�&rkV��eA��VV�4��ʬ	tSEB�J1�0�Z0���{5ܻ��KL�Ҡ =V��	t��i�.d,�M<���(�7��J�����y�I��g�ELJ�@m�r�(�5P�Ym���ݹ���]��5�9��s/�����|Vڬ�P�G)�����e�k�m�ZA��6�����l�"������mNOF?	�$�7�M�3n���z���e{�4o�zm-9�b6����D�0�ޝ�Q���X�bT�P7*7]p}����&�}�:i@_��?��hY��������!���`g?|V�`��#.;�K>�i�T����G2TE}�^�Ca��~���®���t��T3��)�]��e0�����{�f���>�w��3?�+VG�.�Dt����u��b�՗%�[I���L�;(�Q�0J*0�dD	�*p���k܏�@[��z���UL�����L���+��p�d������Ԋ�":��x���3�uݰ�S�@��G�����N��"6�,�6��>�(ؘ%����	�,V����?���I���OA��O���z�ɖ(���3<6X�[�]WbMqsT�dũv	�d{_B��/��b��ׂ;�o�w�f֥D+�m�A�c4���*XWfl���܈�S�+�����������|��XƱ�䐱��TY����pW�J�F#Nԫb�yp��a���@�,�������]����u_��]���mX��G��;��:��k���o���0��3�AZ�c��m�B;�����?6�+�ziӝ�on�xµ�ؙ�p���F��R�$΍=w���z����Qt``H$��?��n��d��HmV�{��V���=���?�h�B��p����|�^k���n�ݔ�·a� ������߃r���Ŗ�m[�ЄN��Ne��Tt,�g6��8��o�N{�ZTJ���nhYx�z���[�~!�^��v��DbQ������/�[�������-K�)�˱i���&'�-I��\q]vҷby��HV4{���H]�\<��/�e��q/�?xV-�b��J�≲�ꓣ�ʺ?��FN��S94�!�Q-�]Vȗ��OR�0�+��K��c�$կ�wM��G-��{!���k���EO]�+%���;e��q�f�����+/lz֮2����G$-�W�	����Y$π�'�]�5eN�c�:�ך bD�cR�]ɋMk��u�ߐ��_�9Q@�X�[#޾�kKq=�Z6k�Q@��ߕ�C����A�u�6Z��3e��$�*��Bo֯?¹8�~����X�o��kw�q^(���1��$<�{�RN����àȐ5��`W�T!�G�����.���]9|��6�☇�,��Zk����NB�#�����ý6�n(���?���mcQ)�����u@r�&����5�L��!$�Q�+$cC�N�*�NA�V*�gߒ��i�����ۦi��I�%ַ�l �3G����\pV�OY9�Ӵ��P�8>������T{���q�qv�5�R��`EN��t́���+�a����%�@�"$T�<<�7*�Ź��<���M�������.)�3?��zd09��k��\_�E�w�f�a�j�*�� G�B����߱Ub�i;/���i��L/
�q���<�Oq�4�k�Qޥ�<�ә�}��
���i�1��v��s��~h��gql��e������6��P���[��Ν�'t1OS[j��"�t�8��E���e
�)�ߏ�b��l5��g�2h��pZ�pt8-���-[3� Q�#)���6<��3��C )��?`����a�����ۢ���ެI��/�����w����%�;�M�7�?��~[]�(��deeAu,ޙ�D�>�y���u��i����~�~V��=���<��gpJ�4M�1�SG���e�ﱞE�n�5=_�|����V�`B��p�j�V��~ D���?|���z�ԛ��2�!���	+��Z�5ޙ������1�A�$+ �2�)��*���4&-$B������������g�8���2l^�HBe=�T~����%�草��{��M�
g�����g�g!���!|O}����wz�'n��;�y����ȣO�����ץ��*uY��V���'����~M��4E��N.�R_��w�Y����/>2�����S��Y�\r���J�>no4J"F�]���J��|_]��@�P5J�5�ۭ�Z~5�w���O�1��Н}���s|��Bto���ZQ��!�GJ����� ��oN��G��@�t�y�d}��(�u,��0Of!����5\���m�ehL�Eh~��|�(	�c�?����pT@�P8�i�K�ؐ��x=�c[�4��R:�Ǡ�n��S����˯#�ł*��qW9-G��r���г�
a)�H������iL[���۝�t;������F�Aͳ�@����r4��i>NT����4r��W3��B�GHx�%���W���(�b8`��u���L�'u���a���x�[�ߝ#C� ��"j��\��I�q��HE�\�qQl���-.JD���� �\o\0D���@Ž� �:�����	����
a�e �)��mP����&�g�Բ.�3>�<�0�
U'	��wu����Bd��pM$[8G�'i�9��S�ض&`��H�iu�
�/c�έ��2ʑ�_��R�Y�#\��\p�6��!���cq��S�V	�=��b%-tRF8u%NCH7�dl\�k�2��j�V���)_�&+_d/d���<;�W�wFgU��Ȧ�.��bj��{���$�_�ځE���&�-�Y�G�@ �~ihY �AJJ43Oc�G��� �?�"枽��t�c�Y[&���І�]'ן��$��
�k��iU���)�M�fl`���,�"����8�|�"d�Х��|��
{�gt�XZ*�D�����6���x��aq+��0�L�_�Dyg!(��VX1إ�(��C����a�4��a2���X� ` �c\���J��;&�/벟��G�&P��/���+�8�ehhGń57N�R��FT���7��
��9�d�TbM���3�[-�A��M6q@�Ȃ���Z���x�5tै8W	G�D���O�����j<m`�(3��Bz�1)¦�ܛ�H憢�0�m)ur�-��ǻ�ڶ��c���\q����߹���>@4�S��#��V�FR�0^z
����!k��p����ă`�rC�	��َj��4���9��XqX\�k�a]E�Ĝ���m�Ќ~���EiQ����<HPh܊��>\���r$��x1���oh9@ζCbmy�����k�^�я�E�1߅��p�K"�X�ݽ�Մ�?:�&$�����İ}�{�c S$Ϣx��vh��-��c�g���s�K�w�,�i���4Zy��v8��Z&�*|+����Yh�r꼹�x��GWC���b�IEO�!���&���d�e�v.��k�,�v��Z(9i��/��81������U������H���$i$�:n�'gsCѳ����J�:qH<�Gnbɍ�dh�o$ן7.���z��Wi�,�؝�0���Ӳ;+��F[��Gu	���P�@Ul[���~��l .L���[)�n�A�dɞ�T�KU�p����4��X���F��#E��d���d�_��~�:���[ݓ�I�*������0����M�ψ�"_�����P���T������`��GQ��xk�$nrE�o�4�I��^����So�*�����*���2�[4┐>:@��������w?�e��� ����79(�1>�[���������C��V>,}XR�]����M�)X��0��lG�����57��&5r�=��iqv0j=����	�7�}A�oe��))���"������"�[Q��frB���뙦ఙ���9�,pjB��Z6��ޣ?���̙B����;T������ߊj�v,#�1!LW���Z�>�I��Ԭn��W�� s�N������^Lp	�;�.	���!��'��K��E�$q\��
;G��� �/>�J���d��P:���!Ų�*x�������ٓv۩%�
��y��X8[Y:_�4R�I4!�5�sR�ϝt��1���a7��e��tS�����w�$�{�5&�vi_�֪OI�\á��_�ٻiSt
���<;��^'H�h��hJ%Р��	��S��bΨ��5�L0�n^�Z�[U0��V�?u�"ܾ(B�a�,l�����^l4sgC�dxOw6�Yn��YQ�d���[��������<�;���u2�*���lyo���n�JE>�0��锖���=T��ԭ6��Y_]UCN�E�r��z0R�_h#,�����C�%��kT\�ON!`�(w{�)wyJ�j�I��i���{� �BSl��S&KUO���̰��㘹vy���NCnHr������_[L��5���G�%��g�SII(1��Ie�E��\F8���@!g'�b��*܊��4�$-�?H�5�����������p&&
N���Q��+�854T��R�7;Y˭U����qZ�Q���k��pq�R+��[�v��\�����9��M����t� �{9]�ɉ���ǅ�9���\z0���ٗ�)SgOa>[jb6!�q̦�ˌ�л�M4h�K�=�O�j�0�TR�C4�sz?v3� ��r��u����e���[��Ʒg���r���b+�����䲲ݭ�]w�_tU��Vb�C�Nn)xi2�p��̧߰���LHx�w�����p8�Pr��m���!��m{�7�ȳ�i$fـ!�m]zBb��6��f[�Q��Z�����[��*Ds���>9�������w�=���u6'5J��_�!\�S���y�2����r~��0 w���t`�b�O+��l�Z��d��KG�� ���i�o��~P�"ժ%۪�#��u湕�����
�sdV����P�,�����.�����1���KJa���ȶ��O"f}5ָ���sl֕�r�I�� �'�����B�Ov��R%cF�ӡ<4=�c�6t��/N�b~��*땎ҖBUg�q�d����m}4A��+�Z��q�]|���5�qZ��|��i�#�R�oĸ��8�[�q��w�E���?�a!��5d�%:ԩ$k���*��*F�U�4����#/�w���Hu�
�b:�����U��u���X �<�rx��A0����"~���2KJ��]ؽ�pOj�&D���:97�д�(���+SΌ��ﱂ���RkD�W�5�����{�$��i4*5K˾�/���m3��Ep`[B"�t���må�s�5�d�
KIOrK��;��U]��h7Qrܑ��hzq��J�Ҳ`Y�m�F*@]ױڍ�+�u���y"�$*��o�{1q$�I�\��A�ÔTZ�o�E�3̵��ҢE�/?��T��~ZC�\�i"E�ɫϸ����H��ni�IJN�����)�������T~�Ϭj�\z���re��}���?<���
�+\	SʴA��ѧcS���P{��ߧ��Z��\�!�A�hx�<�G���!�6�*�S�]�Ɩ4�E�y�){'�+l�}��Xu:�i����-C�6��|+��NN��e�\^�)�]��d�4��p7����� �t���Х���H;h���ҿ��ir*%��S/q~Q����f��*��5$�=ܑ�z�}�_�F��`Cv��Z�bьp�1N�ޘ��)������k�gwLϪ��c�yi�ư�Jv�sq�U[4�ߒb� y�z<1��*HT5�~��h�����J��
�U!SL�JqwgJ+<�΅�XB[�~�8���M����lq�NM,8�75�1f����	��Wqb\ݨΗ�{T��E�5�(?ɂ�7�#�uu����Ֆ��5�跲B�x՗Wa�ZZn��L0�]P��Z�st�X�-˸�d(v�n��ٯ��'c��Ψ�/@|��Bt�\$����3�#��[�*�9�[9��9DG2���K���Ow-��pȗΈ���o��?��i���p9�xǚ=�;�0dD���_�f?s�Xm4ѱ��ϛ�����V��^Y�c�DM�|�ȁ�\�ɭV��Q��;�ta�mͿ��V�}3-Ѻ����5��J�c�^��l=v�,���]���}탂kp�Ѣ5��|؇��F1�y��e2V���s��.;���㊍�`�m�S�䉐��)7��?�����Ζ�wN�FjO2,��77��{��)�E\�MEv��<����-���!�C��n=�͌�Wqk��6`���t�j^�Y�KG��iv�ewr���-�D���١hU|�+[?	�?�k��Z�Y�o[ݷ��$S��Ù�sq��v��u퐿�Fi���
=rZ�k����y�d�]�ݜUe~��>Df��	�����e]S[���PSg�ͦ�"��]+c��:�� ��Х:�h��#��3�Đ`��R��Q��^��23�f}�ό�֤�s�����,��Se����`QL�w崎L�)�𽲒���	��c�v��A�X���ɳ����뿖�K�3�@F?O�*J�<-m7%���1�7╬�� #�AM�
F(�W��YJ�}=��ܺ��g�y�5\K��Y����}?�������%�r�����]���=e���V'�?� Z�>�l�er#R��<6��p���8"�;�ph��e�D"�I��<ء�����)�Z����U�����-��ѓ1�~$e���e>��b�_��.�RI�JLRO����v��4F�(��5k;R��r�u���[�����w�I�OQ�DQ���ֻks~lq�G�������$�� PY1"U��S�{���D��nrT�����z:�����	��p��#��O7F��>sF�ԻQ��ub�7�.Ga�U<��GN�šm��3���GS�O����q�X4����'�J˶^�A0�t��y���%��@�h��w�Ϧ0:��1`i����C�e�#���v�J�P7mCެ�C��:��|�N�@J��������fB{HH��Q*�@L*a�����Q��jGxa}>ϩd���{�!�F��z�^g��A��1�1v,@�oT�G+��
k� :v]�'$�k�#�=�KWm��K��7��ӷU�s���;��2']������f�����U(/p�l=�C��9�¢�s6���(�<}p���m�[��[���H����R�3$}�f3ٴYSh^�p@ױ�6�y���1�j:f��-lk�:4��1�0�/�b�O��ei��y�L�f8�E�U�ހdy���m�UX�PG�R)N�6C��:�Y�3J׃���.��Z���5.�|�n�ν����>Y�mm�_sbӟ��~r���_X,b�EV����]��Z���IikdeNس�v�:fiae�_�����0;��)߄�Zؾ��Hp�jb�j]�,����Ĕ���.���Š��e�
��q�l�Y.L9�b�J�9�h&X��� u�-���|�ޣ�:-ټ�X��%H��4�����Nf�gġ��r<оԪF��$�]����p �:?,4�����6ͱ�-��J-���V�W��~�}�ۦ��K��g�,*C�Q���s�L�\�	ic)��6 +6hg�Խ��U�#���ԑ��ؙފpQ���l8qƪ����RSP�jhX����䌒��d�"�{��c��^�mPl�(9����F����:�c�b�H�8ֽ�\�)�?��J�#��{������ku�3+?���ٵgހ8'�{hd���D(�k��s��;���ʧ�$KJ�.�tk2\D�$ۈ@��4$�����<�)4�ґcRS ,�������O�YQ�	Ѧn?9>B�� M�o�Enm�RX�zM3�4�o��t8ݰF��7:s��1��B����T�Zcz�Ò3��|;G�6��!�"����ƀ�U�F��=ٝiq.P+X��Ob��,�4fߌR���b�0L6�Y�dDYo����l�P���������D�Ӻs���u�2A2����kh�"��"5��i6&��wr�����7`/0�a���r� �����o9�6x����c���H7gī�z\�g������V�U��]d4t:����퀠�.�];g	���b�2��Rm.{Ƨ1�AS<�J��naٕ��^ G��O�oE_`����J��̼���ͽ*n�&��j�>�;�����U�!hf��p��9G'��,\�p�p�Wު�Dmʤy�G64��vp������_�YJeE�նf��#Fфդii���^�O��G�bZ������dyRe�������!:Z��;��R���P��v�@�-C�lظ�9��7C�W�_fZ�3ްg�ا��Q'q4"�s�R�Sb��9ՇPrc����w,�+ؽ��v�L���c�����,r	7-MA̻t�p]�?y�F4�Yn�h'P�1�4wڤ��5{l�e���d�p�J�_�m������Mc8Oڃc\ˮ�7y�df[���<+���/���bn%x�w�� 5{�� Q�K.�N(�Js_Թ�P�G d�E,�ױT^���.��N�"�l�bW�h[���l�v�����ɴ���^ �C'��~m�gq!bHa�"�;ZL-ˋ��EAc���Y��	�_�c-��BEO��5Q@��o[G��0��yEXK�KP�ɼ_�j�kȮ?��ꆢ���  ��$��5������;L>�}��w�u�"�O/y $,�Q��_�p��4B+�Y�,�n�Syκ�������E��u�"<>�!,�~K�m�(tUG�[,����QO�������b,��B�鋓l����+�9����������#հ��&��.C�f�MD`6!(Hpf�^��U߇��<��(۷�⽺��HP~j������T�}V���������Ϋ^��8��<�4�)g��!:��Y++��$�r����q���GX��+��κ҄5��1��j|�M��y��I���),
�^_�\�i�������7��pc���1��!�S�`��@��I�L`N��'��3���YՅ˲�V`���:g����l���u�	 4��3�������t$&���t�ˇvB����G{+�U�
b������� 3��F�5�/�;��yu�.+�r\v��ۃaY�W�%;2���ޜX���z�/K���,)�(^��5�?��Wx��f<+��Y�Y����X��}g���Y�cb��u;�J]_�`�5���v����O���S!�<ʄ�%�幘职Kڃ0�oU��W�82d�O��K����0����5�%���0��Uȩ���9�>]^W.����f!�w���K�c�}UBF�=�omXx�vN5�6u4�
����:] �#�3�MY�]��:S��_��n삶�}_�v��&��f��D��o�c���P�v|�8�21��͜ƌ���i�̓2�ܬ�J&
�������jM��_ș�xM��:�/��PԽ���j��nG6[��: ;JN�⋲LgB6�\~P�/���JgNk�n7{ ��>� $-*���_��M�qHɿ�H�L0�6`�]/�N�Q�u)�C� ��/�EmSO����U/�sBJ͍�8U��|�/�����%�vnwEuaݮcz�VZCJ�v�w	�n�x@�L��ɪ �-�����j���y�&w��r�рs�����cCo~���\7D�#UꝤ��_���l)���.������/W����B���:p�<���;_����'���<��N�}���q����eqs���ɐB���ڳ�ԛ��n$�h�^�`�kIa�FЬDx�[���aHK���o1�"��d̫�H��\�w6\0�PZ]V����?s÷';���i�6��ˊ!z�Y�fjIgw��x�M*�$v��i���G�����ͥ�AH�ۢ-���/^V��&��&�k)���� �,+3�}�1��a2�xV0Wһ,�;S�tF!	��N����7<|Zs̍U.��偤��� x;t��4e�n� +qW�H���}�v��[Q^َUdHo�$�vV���=�`c�Ƌ����
���<p�/����Z�x$�~C��h�8o�ͽ� z�]��tA���5�K��+�`���Z��+�c�ҋ��h�!�Zt����+�UoJ+7�׀���D��g�GS��l6�V�����>Qg�Q!�>}����|�,q�=�f�{]�.,���8R}K6�P��8���]d���ڛkZ���G�{��x�ۺ�UU�nkծ��ڻF�X��c�Vk��bS3b����jD�Ď;Fl�������8�\��:�z���{7��7����8+"q�f�&�RK�be�VH&��)�z����sKi�ƃ�\�qA�7e�)�j���?�p%+Q��Z�B�����	���39D*P�5kt���z%��E��4z4.82���쾝m�fO��k- ,�ly�k~��WY����:��SԘ�p��]~9pb�L�8��á��&�^5��5L��RV]�ɸ��%h~n�G�S�8j��c�K�C&� s�V=t��@qw��)~������J�u��R�*w���Zy��pZ��>���J�˫u3���7ii���O����|�)��a�[?1I�F.Ӹ�l�C��z�߰'ƣ$�����-��r8�8�Y�м���X��Ǉ�� � ���񙕵��e���?_w����A�ޝp�"~��$.�[�C;�T�i�R��^2'uo�5C��KW��g�-��\j0��8ޘ!��7�#�8+S��h~llFfW�=��9�%���"�r�~���'=�X�og֦��!)CvZGIN�ɊC�Κdr`9�2�r�?�VAI��V��F�:_��s�M�W,��]�6��"�fN�PM��:s���W��ѕ��:P���S�"ta���!>�y=^K]�S:�KJ��ư���>�ڐZ�� u�@�El�A�k�#�j�������Ʒ
D���\w�f�U`���V����;��(@KO�=�L���EmQ/T��u�!��ˈyK4پql�x�u�§Hic[�.=���J!��ܚ-�&��dv\y�c�����3��%B;F~A��ps���瀙���b���
���_T�lb�(X˗��7m�P�0�o�� ��f�����K�Qw_����7���":d@;B��7o2���Sjc���?�ۂ1[�A��g�ʋ�O�D������wH��[g�7�R�^'��_S�y�p%e�?��bu�(��?�?)�e���V��i8��������ؐ���/'c|�K�T���M�~���]%�co��)��Òy4r�\�E���u#�:���ɽ��=����$�9���La�)|�G�fgܕwc�uM���ׄ����`Q��+���X�s�
( 8J�(s.�	A�~O�,��������O!��3��5E2:����Jv|w��������QAG�V�F�4v���TP�G�sw!J�U${3�?ޖ�C�h���
��`Ym��H�yា��</��zugo�֌�Zt��aC�B_�eښX���*�ݣA�hx�˦ ��_&�[a2��vwl�59=Ĳ�?�'�ޠ��Q�W��8�i<eo�CA��돞�W2��jx� )@^����F�)?4�-{��=�"����>2Eܙ�S��#os�ȳNP�(�OY���n��B��UD"���m��J�����z=<�X��:��i�o�������t=�:B����1<l�:�æn�ɆY�6&zrd3���C_��J4be1�_�qI��H����QcT�o}��NtT���/�_�C��Eo��m�������T����^YF�^�]q�wA����i>P<Qw����SL�n����d��27w��WeRfx����k����V"�>G�wJ�����O��_3(_ ���5�Ŕ�o����o��8����M�+U����B����� +�|_��w�!���	�3���t�dU;���V2�S6x�\7��Z���a�(�2�kKռ�M�N�PL,��3��3���<��i� �_"��[��^6�/P�O��1T����I���&;~����%����������K�~0��!�~��@���G<C'@2������P��E�C$´�,����4����}i����N��OFZE4y���&R\`9߿��5��B�_�ˤ�5��
����v$�Q"S+��M�_:eh�e��1}ϠkK��ĘC��a�l,�\�������lFY�훶rc�+�*�>鰅�5��>��
�&�����#��T^B�N��T�:oW�.*�t�C�겹�,��.9��v�w�Q&�s�.Yӭ̍��`p�$~�4����d��+�����qD��l����r�3�m�w�h��C-��Z6��O��x���6��_��N��L4�Z���`#U�Z�^L~�{g�K�����l��W\{L�h�{�k�g_��<Ϯ.K&Л�`u��2LW{��5|�$/�"�<!�9�ڭ����%��~n��\۷��6�n��@�;�??Ә���������y��-�JաUC�lj'���r���d��u&�Ē���V��<�����j^��J>:��[�sש:fV�� R�����JL�LW��&�����Dr�B:sg��+h`%X�=��8NҖ��m��E:��^����#D�;N��낶;R�W��b
�j�4�QԌ�>���^�c0Fxm��`~�5{��{����B���{��M^v��"�A���}�W�f�^��K��&�ನlO~1��t���ꈥ�w����:����A�y#�Uk>/���t�w����\�L-[�`�yS��i��Y�\�WU�:Wj~�˼\�����~	)�O	�!N�;Is���Ʒ�����f��q�nl8x|^	�d���u��z�r��b���V@���@���ϻNi�#эE��)ՠ�t�	W�m���r>��Ն����Î(��ȃ�w:i�Yh����+�\r�Mm��I��?ɢ�1wݐP?\�W�# �XW�j:�!Z%�!�o���O���J��.$��%$���F�S����$�����*����B`+���l;�
o4�;1�2�g��Jl�j�i&�r��G��aްw��P���0[�j��<�'Ә��a%l@��l��ov��3��OP�u�����w�i��R�"%�"�]6I��vA!�w5%�(rFD܅��/%k��zۯ�ww�}C2k?�K-��!q�Z����_-s͕��f%]%�@1�Aێ����ë������E_r�M�&�I�(����r0����|�!MY����k�6��TO�n#?��wh\�id����(0kIo��EV2h���ŋ�ސx5M|�=|f].�]�
-�/�@ݗ��������:H��� {� ��"��9�'���V�/��gʺ�]580�����O��ڊ�[�p��XOŎh+����͖9��*��VZ�勪��Ҹ����^�m2j��o���d$���A��N�,��H��R�ˤ���6����Ǣ	t(�Mՙ堀�	P`j3TF�_��qjkB�ҭb��I������C9ϸB��\�*�zĺ+��w!��e\-$d�1G��3��C�{[���.E#ρ a"�k���Nrs���_Cο��d������MA 0	��xɃ��z~B7�e`��hn���@��P~̇o2OƧ!!��MĨ��a��VfL�;��V�Y�0u��%��
h�-���<���8����F:c�(J�0Ҡ�f�~"&�U� ��F�.r2�z�'Z���=#k�HuG�ߝ܋�߮.�?&!���`˾z�e���DQ12)߯��g���h��UP)<�1�Gא��DvP`A	��n�m�aK�Ѿ���i���[m@_:`���Kc6$���z�Aͽ�\\�w?�B�uȻ�������� ���3��u����~� 
�_O����ڛ��CJ���m�;�'�-Q��=��L��Q�y���)=6���e$���+��LyT^�W��Xu��G[�"R����Vq`�:��Lп��[h��ɗ.UU6T=�G�h�@�:������+Xl���W]��#6y~#�������U�\wst(�>��g\I����]9KӀ��!�T�ic�$�&j��XR�2"����������W���� 7�(Z��J�A{h��4�M[�_����;�}y��t��6h��
���.4�o�f�h "[�)/Z�O�
�X@MY6b�ꠀG�ܴ��d	���C�LCm���5�wF퉳�/��+���x���{�3�Ӏ��]6�-���Q�V���̉3C�OQCv��%�!6�$�܍�]�͢ڣ4�.Ej�;�	���e�	�N�uݹ�t�3m�*���Ľ�Ϭ���l�K���!\�П�rE��w�N-fpl��ش{����N��
wk���܌iU�<#��<Y>�����(phץ�㏺�����Upr�U��;���S
o�ec>^
�X�;�7$+kk}z
�w��*���Yk��Ȼ6g[��W��ү�"0�ƍ׫`���5԰a�nx��45���jV}�T�{@lء�$`���ze%�ޣ��I�T�z�
����g]�<d�䛽����i�|��P���g_�<��w��'��q+���m��| � ��$i@���)#��"��c�Os1&h%������%����%����1��������������hcxX�u�Q���ya�wfeM��F7����4�Z��f�wO�Ջ��<��dĝk��N�,����l=��,r߫���|U׬�eȒx�x��kkV���D����0p�×��1�	q�x@4C1�9�{{!O}�yq��i���W��R��Un�)��16[���2Jۋ�*�"�/p�-`[�Fih�V�r�4�����|��J9E���4����z�x�bsvi����3߻���@F�l���6�**�}����e�S�<��$�rspI]���bK�qjm�4��|����g��u[��(�x��z1���f,u�ˠ:���(��*�.��!U#k�s�=y���B�4���DJ"��'�"ɚ'Ś�Mr�,7-�h�Y��ν��(~E�5��á��Ĝ����V��c�2(����L_\��Le�Ȩ4��r�=���H/�w�Wd��=uQ���xq�5��S�8�xtj|l���o��_��y�[U#\ 0KaG�!> ���;�K9o�D���l��%?F����R�D�gc�,�&���3:�?��%p�]5�o���K�}�d����F~>��[O��>�����>���4&�Li�S!AD��v��V���V9ŗd� ��%��_�rQKI
�Y��H ��ޤ�1�> �K
�d�s��Thc��]6���C;C���k5��D#���Y7X�:�w�N���;.�^�'9QD�!Ыh���	~%_<���5۳J�x�e0%_�P�K�f����bg��b�l���w�m�O&�ԅOH�;ܯ���-p}1����?`�ף )��rv�a�+:�O±R�r���=�A��՘Ej�!��<�Lyp`7�d���>�~bb��3�dQ�-�:b'183�3�?��L��!��np�JO#o�`|z����ڕghŌ��e����.p��T�V��:;�F2�G�J}aj�����!�
�jt�������w�[eH
"�J�Ƃ�pr�qzA�筀]�/KT_i(�������\���Nb+?BM����d����;\��&��l�N}Xb�}�����q	�}$)����o��+ƱY��}�n�x�L��IqK�TҐ��-� m�[��C�-���I��!'H� �}�p�>sk��Ϸ ;�v���}#�i����׏�f�U&᱕0�P�4���v�����6�"ƳL����Q;��_�rk���' ���T����'�����+�ոp���O�;�;X����#�'Q�^n�NJ{�;�����3r%�S� �/�����+}gEԖw�z�����!r�]Dڨ��{3��ɖ��k��ɰ�lC��i8������a�j*� �-�t_%X��ɨ��������)EF�ÁzZ��M�'�[���50i�M��5&1���|���~���C��8����i������8|�"ē�8�}���Mtb�?goʾ譩�}��hN�]�Ҷ�$$A�!�B{*Ӌ��r�:�CvN�!��"=�(w��X�������~2: k��^̯k�$����gX��ڃ��H�����I�r��|H�z�LM+���ޚ��K@�z'�h/����F�����mJ#�F�l��1����^ O�U��iK����!�c��L��}b�z�AZ�_�g]���^��@�ROlA ��U)Uw��K��
-3%�P��\����,���Z6�Zx�����d����$��=�QW�mz�(b�����~*%�Q���	(�6���^ʩ�xB��h�mS�����Ι�q<3xk56���]yX�ld�˼�FSe#�M���j��v��:S&$�9Z���W;b�}���.E�~�滚�d�l�}�MM�������3��J�ҩ_�{�-����[v����d�f�þ��I��~۩��5՟��[���a�R�9�\��g@�^~:�M.�n�*����aC�e��ŧ��ؔ�8ʄ��E�T'�]sd1 ��G�~#���2,X������X�,�g�������<���۲�^�l��K�BH({�a�x�T���W��eۂ�d��Z��<���n�\����kg�^��G-I:�=�|V�8���,u������Cr�,-���hy�$��~o�XV�B���O���e����X�:�� ���id�D?Rt)wT��w���R����<��@I��V�������ӑ���B_�%�ޮ	���!�bM\⫼	[ĥ��0h��(Y�?��bq����1ܶX)���F���w��v`1Os^�YƑ��I��W��j��sH_�ǆ�-�&&���|�0��r�s��B�
�����R�_�v�HIR�bJ:�Lx�\�E!�>�V����+�F���m����4��]#Jv�����mΙ�n_��#���}��c8��R �2����+��7���c`��,f�$
�D���y��G6o7Ófg;(y+�]���R56xo�t�'�#����G�;�����kv
���&�5lab�=���$�h����?��[`9!)���0�ݟ��^����|��I~��l�N�7��5vy]�~�����t��s�	����:O�5�a}����f��ݑ�N�6y�n��W�+�,[G�\�[�j��iɦC�l����^�&��B�714sYkH�I�+��:ՠ$k��Ӿ!�����@�}ӡ��x�h#{r����5>���?x�%�-C:u��/W�:��D�z<�y�E�l3^����+b�%��N]�=�V)�)�����e	`��X�����6�l4�o��΀ݍL�M�=:4���ԇb+��$�)�"{�R$ҋY
'N	J0nѫ�����8�����Wo(U�!�9�rb�.�v������"��|˶�Ŝ����>]Z����_bb�Q)����-��K0��eM�������kh�� �W;5�cNyƚ�]��u|�ͻ�ƃh��\,7�����k}/bW<�}�XiU�3��҃m?5���Q�1�Gs�7-�Gd�όmԙ%𝐮*U��v�>g1c�v��+&�0�̢ո2��}+{�kڶ���l�xsms�%Ls&�?N}o�"�?�i�<��k	��NΞ{��&6f��c�Z�;�UE����~O�+��_A�@Goul��@[;e%�I��v�cŸ���v�C2rF�F�Iܦ*j�����'��Q{	-�^�/���`@����S-����o�~UC� ��
�f��/J�Ț�b��6�[\ٻ��1#DE◐nT"z����#��D���������M�Hѥ�Q�nj�g�hs	ox��e�:���Q� ���I�f�d8rC����l�q/���:W�ϬY�̚Y����?!!rk�Lp�ީ�F��V�@<�xz��"�^rȉ��&#���LcRc�X0}x���PЬj�jؖ��R��7�F�� s�EO���Y��R"c���*j��2��H��jU;�FF���c��H>�}�Af��#�3��f�E���GB �B���E�����t)࿗��.rlhڭF���==�Y�ig����؈�N�Z5����|6�����@���v�᥮��@[�\\�]=����lzP?e�p������o)f.�8�*#5^�N��X�P��&βL7���( -c3,�hvu�XR��	�Ü�6���k�H�ιj�u���M�^e��[��n�'�������7,�ALar^�\|7$��0�BT�5�>(��͊q,���	����,?�+�=A0{>�I���^c�'���&��kSۢ1���E�PQV@{X��1"5��@�.wK;��A���)W9��j�Uwn�ec3G��I�0ZI�2���R��". �f�/���u��⯂��hGm ��Ю�%O�%s�&D|���H��h���%أ�nz���O��L�Gz]Ns�56>�/[//Tru'�Q�Ǝ��~�<UE��i�	ˮr�Xg��ۆ�u�iy�nC%����,񐗿Q V9c�xC��[?�$l��Q�S�)�Z��uY�~]�5}���9��Ѯ���k���&�ejam�k&|���Ӵ�F@��ǹSpy��pQ��߳��,�3(7+*}|���0��M}-�&�#T0��I_�f=�(A�����*�(�)�k�Ix���|}`%�Q�#�'m\_��=���78;�o��B��.�7	��)��|y�/ĚqȗTu�k�~O��B��U�f�D�Cz"�k=�!��ZLu��U�<��^(�P1��ީCh�p�fɱ�c�a�hd��lٷ>�Χ��D$B��Z#�ַ\�HTn�K�&?�`�ʨ�(%��jb<�v/�Ht���3J�DE ���!��8��G�+�_ګ�R�U�ܫH8�3ߓ?��������r|�;�IZ�۲2��`{W3�U�yJ7��Ju�x��k��:�]�xY�JD���lJa��{Q�������'�h�����B+1�k��xa����y(����"��i�;OMME�n���"S��D�b���1����#h�,j4���/���d�klپ6pC�B�O�/:ti�&6�E����U4���{CsC�����}�2_�see-��&B3.��!w̫��	�����~5V[�\�ߐ�̋A��^��wFE�Uhj�/Iu2��&C�]y���r\j����1�:k�:ѥp^>4����F�N�J"��.P�I>�~��r�,�1�;W�.�������)�>`���#�i>�/�>�W�5���6�s����ʏ�y�I޾�P��я?ï
�g��Aa':e�����OL ����������ƞd !`�H��hz0,6"�;���j�H������+.u�ha9 ��ذk@dU�����˯B�^�N���sZ�PF������䢛'/�RQ���-]�欯��E3^^���R�����r	�i��l�=;w��	���ؙ��X��K����I��ESė�ŘŔ/꧕m���p�
������pfn�Wl�����sN���<\�#�H���T�,RSմ@#?-A�������gxD�d��%��q�7$�GH�G�!BcF�a-�~1}-ݻ�\Bgѕf���t!�gG�ot��5�����rl����5E��*O��>���2a�C��4��..N�i��b�����������P�����؃M�2g{�����3D��\�����Mq�h5���a��1琫F�v����1�O\Hw<�xq�?g˾�.�E<�+�b�ӚI���~�x��!�,m�N�Tc�i0�������"�+��w8�?Ug�m�ϯ�"4�?�T�`W�n�RU�8L�n�%Gok c~o\��v���O�=����>L8�i���>�3|{�b8��yC�a8���O�s�t��qZ��O3�^�D���8! o��g_��B�7�&����V�*���B������ZI��\�̠��t^Ek ��4f��4,�������)Sۄ	�D�'���{__.X~5T�5��.6&�0Tw��A�څ�x%V�aƯZ�����{�l�$��%�R$�����n�cVu�N%���|��x߷��y.>:Q�l^�p,S�#��d�U��ѹ�cX�៾��7.7Ⱓ� x��]�(����� �z�a���f�WT�~�Q���o+c��ԅ�d����J��ٜ?sf�{��s��I��JK��b��t��o� k�ZtN�/ԇ؍{��޻������w�Pwh��T���5�&�J^�XFt����3��8W��w�]�CXD�+�h�iϏu��[Wߴ������[� w�: �p('b�I������+5s�z,��4��cv�r�kn؆����Is�׫��"n ���Q�����Ria�n�A7��V�w�1���Kއͨ���j�yAa�kY�JTE��=�&����Xw���r���Jo�+{s`;�.�D��ԢG��y���1,�����n��A%r�LPyrhʕ j�ݻn;�8��,�TIH��i��|�\p�{Wɥ1:�K�*C��-� L!��X��8��A�j�p�d�o<���-xqp����e�<��q�OF����_��Z��|%[8�;�#��jC�����~sn��b��h�^�^Ƹl{��n�ں;���@']���~mDbC�g���Vrޤ�<�<4��o9n��CTip���1}��5ё�g����w*�O����B��O����M�o����DX.*�r���˝����:y������ۦ@T~���ݸ|�s<v�̦ˋ~ӻ�u�"pFh ޺��*H8�-���^U����=���o}�����v�,��W�r��o�N��a	��*^x�֘�
::=�2�����g��N�2~�����M�k�b1��4�I�l�>c���WC�Gŵn�;�7O��ŁH�mFԜ�V�X���-�A��cCJ�i� &��I��������qĳ�9�W�:�G����b�H��=y�;�ta����͗����ј�[��-g�"s�;����@4;49�>���V28��nYcN����s:�Y�".�儧�%���p�"��M�к݋�<�F1�;�_
��N0��	LJ}o�G%&W�+3�yŅ�o47�%)�,���D��t�Փz��$�@�<<�� �RG?�I ��QKϣ튪T���wQ������%�L8�@�(ө�@l^̼3��:x���+��X�\04���PJeI�+�T���J�U��'�����)z~�!
=�-�/�M�}����Hr�hl]&�9&ۤ������i�OT[��˱�1��]�	J������},��A/�yKӐ>��\+��p~	�l��C�7B�i�i�B��+]|*�!T�
���SM�4ΨF�����r��� �k�µ(�NI��1y�Is]���y�#4=�UjK-K���#+w�"ͣ�0!�K���L[(�1�oF��t�K^��!{]��vi���T�ُ\_��G5�j��F����7��2���5�X��6����M�[�*W��2��H)>Z�{���wH�$���-��j�����Js�(����餪�G��<p)�%��I&���5�z	���7�t�(M[N��x۝��3��+�8��9u� 䙱�i�L���� ѰL�>1�6��I��O6����R�?���CZ��
�5�Y猖�A�����uQbY�U��b�-��ٜ�w�w����{ot��O�����[#�_JO���K`1�T����=u,+D��3|�֋��V|4��'���e�J��]V2�w��4EW����*��X���J�B��N�Y�4�SX>1�iz��C������Bs�8���T�l	k�4Y���Q�	��b̙����'�cB�mBO�tD3�����6aw��R	��V:����7�)�q9mb(B3�ϻ��E%�/��=����K2(p�k�}�smrAR]�N�I�&8�� �2B_������M���Pѩ��{���P���*x�wnV�p/��o����[�K�@t���7k�;:U&�9HT��GbT:CHI�sW��/>@VӦw}ס'u�#O�W��{�	k��Q��r6W����M@��5c�~I������&{JE����Y�O���DZ�B����f��3�)��¯dQ��q��!��x1�	  yY�s���cq ��=d�p{bdh�mr�.�� �("�����=�ycl^1ͬfH��4���ml�5X�4����p�tЍ�&S����~
w8�\Y���t�a�G���� 0�����7��BC)�����u��Ϊ?����j�㠨ns���F,wBgN-Y���j�5��8Q�w0	�	��&��n���4����L�ˊ����C�=s�4 ��PZ�ʢό���t��>�7v;̲V�C��NRq���E��a+]�l�|4]�y�����Kަ-��?����b�N�ي��/ѫ��-�������تڃFg�W������u=����wV�����D^��GIy?@
��6+yL����Ɇd�J��"G�gcѡ�1q�`f�"�Ku�����ض߇b��
��.���]���*�{gXq���7��t���K#�����Ͷ7-�#6$�tǲ �r�FMF|[��	v����(!{v˸eԔ�`'�?5t**�S�|7��Tk5�=��`�K�t
 QQ�>�����:���OAʥ&�Ӧ�����T~��ra��9%ܫ�W/�o�Gr��'�/�'[��7�M�'�1���jӯ>*�(M3sK�y��¿2:���4_[�o�%��K��qF�XţPS���,�>]���[#�rܓ/$<x� cO	��\��S����Ij�����m��d�'OnI'ռS�5�X�r��e�RBu�5ə�C�[@�5�Se��0m�SE������,f�@�r�
wi���"̌R�0�W������C^�TWqr_�e�ߐ�aV��"�����(�"g�&{w�+<mv��^�R��F���bH?4�d�%�z:-3z-���;;:�F�^/���Z����ţ������)7�ؿl�(�5�?J�Z�m�4�ع5�_�ʜo��gG8�`o)>^��e�Tb(�;eU�D����ڧ���x������ޖ�!\�h�T�_��`��p׏��v��؆]�&ț�G�j��c�F�8� R�Ě��&#cinx%)t�S ]~ �2ۄfC�Zg^�?�nÒ�.��{������Es &�FGT�i�5~��i����1��x��'.��)C�̦�"W��3e��r���_Ӭt��&�M=`�ׂ�s��b�����=\�	8e4t�������4l�d̸��`�~���΅����?q�՝9�~��e���M�ʜ��j_op���!J2=�|Ό�~S��3�F���E��wA��`�@�Q�9�~��]������;L�E���]�l�����w�%��=,��,<�I�����C���Qտl����g�����l�'�"���M�j�����Y�H�{"5���߆2�m��.#}������Ġ�u&n�X�5)�?� �$�e�+�GF!~�2�o}�����9�D���QP&f�fiU+CrP����w��N��c��8��E �B9�	L�o\�d�����;�v�3�p�^wj֓���qTV��(���C����k��������&��g�e�]RNSo����)=��oHؐ���-\_5!�ߺl`�Q���ZS�כH����ݐ�WٓAA���Y�!�q�Cd��G]��%<��9�u��qy�w=e��6�1w(c�Tɵ�Q��>�����ay��b0\-Jb��x�D����ϱ�ԅqpq���dS#���9��O/>p��S��6��fdFH�	����7�Iݡ���nN��Y����"/s��P.���j99���N��m��6�鄢�<4$�tU5,.�y�ܐ����i�LA�E�����N%4�1�8>>3����y�z})��i�,�;���w�,y�`��,hϠ�ֿo�25ͣ�,t`9]�1�EfCƱC�/\5�h� �:�$|�,�\i)M��1R����
bN{._>�/qM�3����&��f���j(�5!���k�E$ݿ!ڕ�E��<��A�S�n{Q��/h�*:�'�^� �{�ɵǊ{I�����ג�x���N����&��T�e�
O�����0��0�C�r����߾՝�1����f�ԍ?�������bu���<�ζ��-�V���~�{Ͽ�p]�����8�a律KS���\���1Cqc���[U�L	����G�ۣ�L�Xݧ�u��cmb�2h(�h�<��M��Мf6q��<jx/�9�g��a�U�-u���㲙����R�,�����ƭ��tg�0���������|�.�0p ofu���w�����G���l<�����DV�,IxZ�$EL������!�79xr�m_m�G,*��luŗ6��z������!ِ�Sǔ��s'W��;�<� ����q����IwP���*o�e�V��q��L��7+��Ut�T�s��{���D�9��ȭm
o��0n �:��s��h�ύ�)OE?�H��/y9��l���ZꖎCN������+@�g��N��oHꑉg�S�v��;Sd>D�0(;�2h�Z²�ސlwT{OAv9�Ĉ��5C�B?\�J����E�ۄ���=��pG�2���H���g\�	�!���(�;o7��$�2X@�ۉ���w���u�W�6��S5nNW�!��fֆ/_����6�bn�º:U��`�Z�����!4��Լȧ�6�$v)�"�Gۜ��e9�˂.u�5S����3��k��j�4o�\I��io�d�GY�{`�&v<��{ʖ�Bs�#S�x�����|`+D�r#gY	�@	�cQ��E�qr��w3R�	�;�¯�sE"��P�ɩl��6H����04�H<�{z��&�I��BV��xՊM�['�'1�l���7`f������+z�p龖�����C����̉�1�ȩN�����㧑�6B���xWf~3y���L��}�h.���0��i1~'���߬��w�'U���37	���9�^�C���Z��W|�W�տu���D�jV�������M�N}�׊�qզ_�$��$c�v�Ѧ����|^��'�$]���;@�Ȕ>���+S%�<���w�_h�5�=���W&|���F�UVk�s<M�\B�����oF����:��z����sxy�M.���\eU�,բؐnK�ֿ�!��-��ӽYKMt��4�B��T��>���d��jQj��U�5e�c���U#.5o�p�+mA�-��)�ַ���"�����7�]��.RW;�Q�.��9�Nl�%�ou؋тyN{n�
-;�j�#��׈ 5�<ѣ)B=���dO�O�{+uT�xI�������幞�|a	o����"g.V_C3�`cubyi%�57$�\&>D=�Ak�S�ۃ<Yg#_Z�Z�U��?	ܾ��9�THIHI����6�$E�׊�lH��r�y��K�:�����β��?�`g-��/�P���P>y��E��Q�v������fC\�ֹ5��0
����pĂ�3��t�j�`��7�'�Ze�B��C�Ͱ��"YK\��a�Jk�Q�q{L�y�CYs����F>��.ty�����q�NF��^EKvO��w�×�k��C�&V��£柪A�1�,�!rm��d�(������tĶ�M
��ڃe���HӜ�ڟ��k�~��-!Σ'|.P��jN+Ș{6�O�Q9vީ��c���|R5�:�T�j-��ׅK�T����̏]w~���������M��M���f�ydQ5�_uV&ء�dHp��.w���G�ٖ�`�=� ��yN�	&���&�o׺�#줎]I���%ʿ��.T��Hms}�P��A�@(��]�XKs`�s)��'� 
��~pC����K���c�ի���?�9��O~Zˠ���*?�f�^Ѥv}YX�R���K&��#��;j�ސT��i��<ڌ'/��h�0:������k�/��Iο���D�*9w�G��i��[ɔ�M3���܊[w�j����:D�,���Q'Qe�VZ�� �TC�ک�y����W��
�����4��g�ʋJ���nHx���`�[ʘF9*����m��%�?���
��H_�S�3���fb�Oc�fӸ%(<��G m+�Xk��؍X�ۓ�-D*9�O��j��a�"0:JhO&QJa�NP�3�-8N��Kd^/E0�α�A��(c�oe��rږ�$�oW�Y�c�b��[����[��=�" R*(
Cw��5t)���(H�PC���H-9#-Cww�����������<�׾�Y��ב��}��&(Öو.�x�ۚW�\ױ[� ���q8;Dۏvr1��t��0�B�sg�
���10�j5)�@�E�U�|/��Ft�C��Q,aF�R��>��V���{YҨ���s�'�3�m`4ڼ�f���e��Y~�R<�g^� qUH��l�c�!��N��k
��>��EN� ��O=d��Q��S�d�u��%xT�_Ǽ�4_Uu�{�{V��݆�j�้��)"��~b�*R�2�E�,�Mwg�?#=6�l���ܟ�I�����7�	lѦ�wn3���_��c�{�h���-h��.j^�����>�"I^h*�(���+�p�8��_���b�E�5���Z���n0q�e��b_T�e{����}gv��G[����� ��]�	x)�[6��r�,�`�����c ���٘�(�=�p|Ւt��mwy���q#te{���d�v��� �K�����[1�1Ņ6�(���E5[w�(-�E���«�'i�~B^tl=��̔N{?�3�/�|Vޠu��4�[�5�a��e3�Ħw��w"����
���Z�,]uB�<U�^"zsד�#2�2�����cq��8eZ\]ۻ���0Cy��\?�fNr�ev��j�\'SR��PNh���+?��ԣ�0<��Y^�g�n4�e�8����� c�v���ni���:��9k�8&�H���
����^=i4�<*|?����1E:��,��	��c�BV�6~�������1�J+Sph�����k;����� �[JA=aNM(}O�r)���~�_lvv�}G�r�-2�f��H'.��oQ��E�;��"����k�g셪�Ԯ!��T��f�����x�7*������PK�+���!�Ño%�� |wƆp4�p$�H9�W�eq�3�����F��ij��L��f���.������1��GVmla�*�g�{a���Gۙ���&k^ҼAN� �t̯10����f��w�$l����8k�(���n?Hqb ¼��6�);q���gP<s�b*���A�9�������*�W�oT�6��a�Ȋ)��G�����˵X���O3�V�;�$�h�)p��u��6��>�e���r�D0�>��0�m�&d��ķvY�e=�}���3���(	�o��?�[]rDn�z*�-5w�{[a��ǲ��AuR�4!8��B��K�{���8�O!�X�]6!dx�0�:����&,j�p�S�9���5��Mk�z��+yow9���$wiM���~Ii��O6V�ۭ�o�������ߗW�h�ퟀ��}��-�a�BG- �k��Hx)je
f�t0a6�P�[��x���[o�8���y95�lw��g"�<���>Q?p 5�<�g�%s�^X����y6��<,��r24[���<\Xׄ[J�m7숶j�hŶY�w�$e�/��RP���
n�W��;s�����T�Q`T�ǊDu�F%�K�Q���L�*�'ɮ�VG��W��<�9��~��QNE�<��%S��~W���`������\>�/旭`��&�vAڔH�������s	���@���?%#�AB��7&�3[�o��C|\r���0s�^y��^�������0�+B��X1g�k�5����Qdc"��%Bb|~�n~��Ҙ	�]�3�}��J�H��l\߁GKq��m=��g����e���Ȟ�U]4c���`Z7�)0&o�[0ѹ.<�������I$?���~��O�<��Rv]7�Wyx3�L0�G��h~�P�����}J��:Yl]�I`����\�*���t��?�o�m)����ɽ���n!}:2%�A.<���;��ˀ�=�fb�;�I����@����ўI�W�	Y�=�����p�V��I��̽�����3�R�:3g��e;��v?�|���� 2��}P1g���ک0�/X�vW!H{h#!�=	��Ϭ�V��؝���B�5C�d�_��L�+�,���k��`O��ӕ�!��#VGp"i8}"w͋�����#����!I5`9�}�����'+8Yǟ����\�R.���>yv[#���=���*.N���Qb �8P-�ōf��5���q)�Yڷ��e��P�"�9����,~�n2��� ��]��o���3�*~��Y_�C�,y)�}/�7�*���L��&�X�v�q~�ҕ��ȑ/��S�d2��f�r�5�L�R�r���k5�4���G(���iõX�7���X8v�jΙ,|LD�s��֖��GդX�8�5��m"�w}}}(ol����|�9��8��WmPk_��C����;���r�@6@	i�6�n�o*�xi:'�G��nt��3[O�t4��.:��]�To�rl�}^%���=^�������M�H��*w�-�>�|��16@%W�달� ���Zb�ƛl'���ͩ|�_4k��vgbH�_�'t��%�.h$��=��b�
�r7��6佰9fO�#�_=�M������'A�*�.��UII��}1���*ɶ���9���H�La�z����dZ��b̥�����^]~������ԩhe����������̳��R��\����2�E�|I	�Y��i}�쿹�ҙ����+n���`b%*�cEڅgm�G0�^�MA�G�D�f��WM�oC
޵u0�RY��G�u�`��I���SQ�VX����٠�(�6�2
v�7:ٿ;�Tv�J<�v�aܢ��~�t�~�pEMfzD��J*<�=���D$��d����E��@]��6�e�~�O׽�
rY޿��<�C9���'�8��l��W!���:��:��Y�l���˲~<����͒��A$[g�Uv��ǰ�IPn�v���/��Ύ�7%���M,ۭ���%��J/�����
��xkʯk�X�g�3��xB=w�&��sK���9m�a���@)�Q?�q?��K�����]�'��½��~W��̞�US�� D��=K�,޼����ྪ{a�Ѳ fv��@���$�k�#.�5�+����N�/��l�%r*\+�.�A�`���
#x)j�~VG0�íUi�#������zBs��~�\�]V���[_8�vT;��a�>H��NY�*rxn�v\��
�e_�2`����WW�>����A�֠g��>Ļ���������u��z�W��z�Ě@��5� �nJ%�����}�km0#ئײַ'��v4�Op���pL�B�U�+��-7�W������с���IgS�b�!�*�������"ٔȵ����J�94���m �>�R��}����ϐ�һ�w��j&P���d�:Z@���.��ȻVj�!jg5+}�VT%<�X���IcS�G�&�o"�~""F�1�D�q�.k�t���b�v�$�)��K��¼A
�J�[�a��O�J���s����:ޏ�9[�=,8[A�vx�x��_/{����(�S�y���4��,7�5��V�6�$�8��s�j�j5��I�ӈ6:����M-�{�8�Q�����7ͱ�eRpb؆�8�8k>�q�<�)�x��#�X���O[�Mz�j�9)W�V�ddroC�^�-[V��b�\G�)��6��0�>��5�y�==�j|GV8�.��6b
"KV��~S<�R?�Z��3�j�[��Va���	��!nIMe �"�V��z�RP�A���k>��	�R��,���j���I���4��p������K����M�7�yL�=��%�y� ����Μ�M"�a�፱hmX�aۈwHh��c��ٕAy�S���ɻv�Dwۉ�|7���ކ�HB;��mE�I���90w�{"�N�)��H�+��w5�����qõ�?��e�TB�OFۇ�u]A1�h߶9��V�]L��!�ww���~���X9/j^�䠢^r}�PE3a���%l9��[v���A˲�{�hV���_��>�C�*�$�^9�:��Sr��j|�L��%�~����ֿ�����F���76s͛� �A��'p\@�����s����|��V!{K�5fL����M�7ժ�C�xm�Ll��Ht2-r�VߛNK��">|љR����ێXAǌ���G��H�`���#����R�V���u�P�1e�`�k�lVd���K�R�����ͧ˱�l�\�j]�rȉ�\�-x�}��<��Y�y��%�f�E����~�P�����Q�|	}R�s0�����so���8��0�ɝ七����CXK@���b��_�b����D�;	���"����m�f��uiii<�����f�d�^��Y=��<�q`T	��z
�}�������1~s�U �?A��>L���y:�N�M��%��;^�A�1�b3l1�Q"��z[Z������Py��6�_��_�d�F{��9<J�<�$�_����´����5����\��O��p� ��[[�R��ъ���B�E���u�p�����#`$��;>^�&��a+y��,�Љ,u��/�;B뭫�.���uҟ?>˙�<Y��F|t�����_�ۍZ��d�����B��sKL�v��O�#�����~��(`W�ֳPn�k�~�����eX�0skSL���xy��Lǉa�R������+��CDjo��&�U$�>��*%e�2
����"DV^��P��X���ueb.��&+��3I��qI�?�p	:�_kٟ�@q9>r]:	��Ѿ�~��10ĿD68T˯Ԩ+�X����.��I�������T^��ղ�$�q�@�bXG����9f���#���ޒxq�+�bQ�n��U�n�k2n����f\T,�+�K�@��Li�WE��*h��Y�U���9�k�7E�^op�u1Q�R��	�ʺ��x)�8(��qd�.��.���k����P�����>Ŋl��Z�<(�27�S���$�J�Ä�EC�qR8fS��#�k������>9�ߏ��s��]�`�U��o4S�o�/�Y�K�VJP�:�)��f{�DT�-��x;]*����JR�G�D�[2���4�LJNɏ���f3;��)���z��+�G��y�U�L������P���>�El�gAj�~T"�@#CV�����J���`�6
~�0:�kH�]qD�AQZ7��[�`$�Q]?Gs�Tv�p�g& w��%{9aN�g�|hg��w��g=:�ߢ��2�M[�& �~a;���-�&ݧ�N��L���^)~\�����(	E0I&��B'��2��:=,�E���v�O��h\�a՗i���/��PB�k�E�@���t��&l=-�_fh�MV��^g�ۇ�2a#�o�N�8ә�;\g����Gk��3�G�_�?��P��ۏ#E�FN#4bg+�.ݨ����h��p�疞g��D��dx��f0E����S�����	�+24B�����D�L��0�CEI��8gN������<\�J�m���G@8j�>��2�c���2imzǉ/a��)��o�or`̩����"Q⌛q��䨱0=���&4����c�4N
��e4��5���1G*�<���z�\��~�(+w3���-Pi�hj-�Qh˩*D�f�z�DcXl����'VEp�|��r��G ���q.���}9�{e枸>*�<e��˧������+˩R�x�׉�NRP��W�N���L0�+�����ۭ���P{AY�[���+�W�9I����ddזU`+�PW=�n�>:��\}�?p6�ZQXU�D��$�A�r.��,� �O"S�<w�2C����4��L��c�ǿ]��'k�t40L��̖,m+�4�@駈<�G �L<��z�)��W����mէO�y�������rU|.�{�[�G�6��UK���ܱ�m�Z�g^V;���"�� ^��C~����"����F����92��$����	R�ʏ���NK{�S|�@S�
}H$[5G�����v�>�������#�B^=.���:	�yѬ����V1.PH���ڟ����ܘ|S6��E��7=g���T߄P�\ul
�(UR���2N��!+�Y�m��ˊ/6:ynsm���9���9�]F��T�,�!���
:|�\��PMN���L���J��8o��0�n����șj �kR�jජ��DYV3��t�E�6��Ũ���b�t��<*PM�I�6�}Va�͗8��l�W������i��>,O�Y���E9���^��-%B����0��:��@�H,���`�G�aL#�ؕ�a$�SJ�L�c��r���fȝ����6�T\�`34�QҳM�=�`m��c��]�߫�S��~عu��ɺaC��O2o�E)@Hb_���$Dm�x�`�z1��N3��V�؞�k�~2�`��t�zb4��n��uD���K��)���B��ƛU'$?\%x�����1k��������3�N+Ɲ[Q�l�أ��"�@��$pb�Ϛ�� ��eD�4˒��<��爩�<����������p,��1er�>A�f;��Xi�7H�:8kGu"�_z�B$�[7�x�f�Rh�����X�J������9X��5�����t	�@Mf�!��F�SV�RZR�ٹZӋ��s?���y��X�h�7�cǘ���7Ց�8*�<�.q�ճ2���0)��uu�"�a��J�To����H�'$�m6\�K�<��8k�';��	�q����d�ͽA�0�^��T��s��2s�^��ޛ�\�p��#�ϿH?o�z�^�bB����:� ov��7���17�I�Yk����_Nq�?��+2)mEU��s������&�z��Քdo��'����ٿ��ΞOa~�P؋��ؕ�+���ϝ޸-FsD{��e3�4�:]bbnJ�<����*�ݏ]7�C{���?���L�:}K:\F�����e7C�B�C�w��76�0]dE:���5W2��5���@��E�U�?�r�5xw�t֦)���	��/�Ǣ?íK�6�R��+����J	[�Il��c�O�=~�{�YiS[,D��\Nb��Q��m��}!���n�pa�ߴ���d-�ח�����T��KK}���V���ﾈ�H�ך'qe�������+�?�L2�G���r��#v�w�!�-"�J������z����:;�vn�~��2fO�2�ܲ6_\�~�㽑�y�YTl�;�P�����?�]M��'f���'f<��	 ����sV~8���v\�w}��ċS�f|<��FbŤ*�4r�oiW�r�5�}ЬSM�x�	���
:���E�J��TՆ�/��֌��9��j?(qH���ΰ�H|G|�I���N�l���˷��#$c�<�S�s�8��FM����۪�uR{�"�	�ܪ[3��y.��1e/��m���~���	L������F�lr�Տ}�ٵf'��Kc�:E1O�R[Z*0NKJ���6%:��I+�>[��n�*B�A���Pm�z�MD�9��T�7�mis5 �ۭ��"�?hٵl��ury'�i�{]o���}�DF/��n_�Eu���a�}?W�G�ؾ�����ÓC!A7^�?��j�Rf5��`�xE;ϟb���:~ƻL��7�3v��8��976�ު��;m�N��%�k��is��eXg�������x5�-;d%�E�
�x�$Nj3��rt�d�iJ�*C���WM��m�vXvG�b?�?��{:���D���y�Y*�1W(}��
�$GL����t�#���r�;zr�F��O�ߓPQY4�d�q/����iBۤ�>L�ۖ��
���4vE�������~tGw���Q�t�`���1CW�c�~�>���YPJ�ߒ|k��"�Y��8u6����{$�����!�ԌY蔴�b���/m��V�4��U���a�����ߟ���)��+p�N<�1��z�oq`���~ȑx���n%(�\#5�fbu-Ft_�����H8Y��x-�=h���ٍ�lOjmW��u�uq�UMg�GדŬ&�4}_[	���-�3��-��Q�醭|�ؾ5#ٍ�f��O�f7�R�ה�1�n����U�Х�O�����,F�LH=��"�L3~4�P�,�l�}��}6\��5��,�}�~���`��=δz��A�0��� ����6��t��2���\U��Y ������w��v�ǞWMY��2|��;��AWKCt��m/6�l#[���c�^g!F�Ue�rX���BXs~�������Z��M_oz��c��.F�5�]^�b�9�M� =�y��&�Rd<-ޯQ�_´>d'6`�.�������6�´c{xs�KR*��Rr�e�q`q l�" �֪�	�K9?S���c|��p�\!�K�Z�,�Љ�ç�.������	�N�����l�D.���=am%#M�����=Cn�r�ŝm=�$�����2�r�A���s���?��ֺ��С�C�V�g�+������;����-S��.η����L-�������Jx{�>�~V��A�h	�Y;�`'Ѩv�@���Dl-&��8����=�x7G-����bZ��2��I9���g�����w�{3��;�gU+a��6�v/Sq��.ʁ߰|���!"��V����h�Nꑽ�n�l���4o �nݝ W��>ʾ�;��IMY�-�M����U7 ɪ���w����~C�����3w�Z��,���r��%Y�FS��L-���5r������N� t1W9t#�OL���� ���H�+��[V��E���3E
+@"а)�5p15V{����b����^�2�=���Zh�]��gn^p܆+�Aa�l���ȽzQi	PK�H�cA2#GM<f?c:SN=�iv��R4�չ5��N��՝U��+�aHu�W�롆����E��Nw��u�����ѧ;]=�izS�3����~���D�c���=jL��pR�=���qy������
���Y$��u�)�*�#f���A��HB�����O{E�<ϵT�eM k�ME��~��5�(.�����ڝ6�-n�jۥVA�k�_���'�rc�r��&����h���hu<���
��14>�x�A�u��:� �rm��2�I�����fd�R��ҀZV���ʠ��T͊��̝�}x+V���~�r�?ѓ~�;LՇ��\�����
e����Py�i�bk$P�6W)��%��A�	��\�(���iU����x9�խO}j�ARi�UvC�g��ȋ�,�m���B���d�p[$o;���v3�� �����<�-�hDܤ4W�����{�ŏ�{̖���Ĝ��f��%�x-����br�;(Lf��s>U��/�#Z��s�=��Nl$�25��`���{,Lѩ4�X#�
�k2�T��U�L��M����6
�;���r��ث�S�x��nP��|��'������O��e���Y�5���ܕY��9�Ȧ�S�����0��F�G�WZd� w��G����̿X�	��""v(����]�I����]lЬ�__���KԳ�#<s���\P�.U�D=�����y���>R|�後�����M�?���E9L�|��}
3ߠ	�w������+)t�1�%r�e�`7�*��=ђ��VQ��gi~�����ks'������Ԍ�EI)�x�b_��tr�≷&F+Xsn>��P��'�� 7t�v�H�}�E��X��?!Jƞ�*��H��.n�b� 2���AɪΪ\oV�"��m32VHy��̎	d���gi6�hc�ϫj�3X�ӳ���ڗ��׊��׍=�����^�{/���|/:"�9V�MAؔ�]bM�59�L�a�;|�F6�Pɧ�&��d	�_��?�}�k��uJ�m�%�P�ꩧ�|B<t�ȫ��V��d��
ng+��OS��q��2���}$�3Fa����A�I��ivT��jt	�h'������_x�-I��ϒ�R0Tm����ϵ*�����6�l�I3m��_�
�Ћ�N,v-a�Sii���TzPT��9��*ϲs���.�8IϹV��N��7r=FJ�i�ԁ�5Y���;���-PU���f[�5(I75�{H�ܣ�R^��`-CѠMW�+��P�'�E�ܽ��gy���S?���:a��9��:�G�B�s���h
/�a��mI|��)��.�ū�:�E�t�*�)���d�zq��R!t�¾��4v�o����7��_T�r� u]��=�:��֯m7wp��ɵ:pn�	���kI��LV�,ƲL�l�A���p�6B�٧�sb	ʃt��!�}�7 ���q�=��sֹVs�璒�5�lLx���.6.�F����ݢ5j%1ݸ���M����u�2�ޢE�,��Ô��y���ƶ��D����D��u���(6 w�&�p� �_�goz�Y�����rQL[*��/���6�0/��>e���-�a�[�c2VG�t��1�e��T,����}��RȽ@���-/+�3uyR��Mou���V,�P\g�P�W�"��1tZ�M$4�ŀ�� >��?�9L���yy��@qV$�o�>�����f���7<P�`�q{�t����Qۋ,N��^?�gq��I�i�E�+�cY�(mW&*^!*�bN�a���x.����Os8�9N�����+s��H\�Z
�4�7�u����Ӥ0^u��@b:V��Em0pTy�/+۬�K��]������s$���_�`o�+G��ڍ~�4.�Y��H�N%�̕"��{i��~�������hc5�o�$�"|a'a6~.��2,�#u��>���%V�9P�x!͒ÂiZ��Y��ֆ��K����|���ث���2�@|�0_l����{/��*0&��).�^�l#�c�7&AV�Q�����3_
�Jdt�ד����q�ȟ(`�"����e�?)[���oكE4� ETG�-���v�����Ӱ5.���XhaZ���r�C��a�;D~t�d��}�֬����v��x]��ҹNV�랉K�]8�6�e��\�t�ǟs	D��f�7��mn(���}�>���Z�����_q��a�6������~����D�Y�ɶ5�u�m�K��#)�,F��9L]�����Tp\lW��".�	��`R��ܮw<l��-bǡΧ���ڧ];b���r���գ�I	��ә�>��u'@q"S8��Y,��v,=����Ilv����ݲcx]�����s��+�N1��_�uͶ��}<Y�z@K������7�֑b�8A���B'��-�0�Qr�5֍�zN|���i��%gj���`� �Ee�*�^�?pQ�۫�l�iz=�� ���52�p�\�g�IO�8�o��7g��{���� ��Y�F;@)��ʮ�:ф��d}f����Xǎ����s��� X
�M�`��>�>..�{X�2���ښ��[c���%:T.a?�dW�����-p.�^��}��~A0p��q��Ӱ���i��Q�_�Z�'�hUk�Y��蘮d�^�m���7��ۜW�qʝ��H���>8���A��C���w��k�YW���v��܍Ĕ'Wף�
�m�
���	ڵ�:C�zt� zΛ�{�DC4SS����h�c��:�)����q��Hdk!k��M��y�g��6'	�lX?Ye%�:ҋZ~��)�V?'���W��b�>�v6�C�M]t�<����@Nj�n�'[�ު|e(2�B$�]<�|U��z���B�"r���j�4�څ�b��Ǽ�mp�d
	>��g�/+W�����};I��XW4��+����5����\�����B�����Z��t/�b�D��MZ����nh�ń���m�,#���^���RrN��(;bVģ���$s��(0(��ڏJ8	X%�n2�ŗ�K���=?`f�����>��i��D�E>��Cq�S����˗/^�p/������
�������܆�^��G�U+Ƶ�R�`�d�� QgЧ�}�{v�#)7�)lb�/x�e��?�\0G��'��&���:�S�8��	�����J�F�I>��&D\��D�8����^<pIN��ߵ�_-�ox����W�g�R�m�d_��B�^\�.w �
ILw��.�UY�4㷤�'���,J����_�������X]�cz;k)�#��M�8a���T��́�N�Ҍ�S�Ӛ�/nd'41b�`ԚyCC��# �w���k!�m����j��P��|�x���5�#/�5G�ف4&S�p���:?}��(%�����l�kq�`�`�������6�󚆀��(m������n���49v��	4�
Tc���d�_����
E����s�[U��ƅ��k�^/��1PC�!�
���؂��.��t��gڰCBϡ���oc���I-��vn��a��ã&D��>�&����J�܁:1�WI�d�4c�&x���bt�j��ׁ��ON�:r��i$I���~t�Ճ�B��A��4�Emo��z$%~�i�jE�ʊ�/�^(���:�x� =�`X��('��r��SL��C����\����D����8��t,6�Y2B ǴE{C�f7�B2�:�,s�D�)�_<�?�Dk�����fx�]�k7ӔKG�yPZb59��x�s�&�<������Џ�!d�C^'���d�)���e��I[n�K{����xUT�*��w�)�;&7��<b��TW�
n� �Z�~#�!��w��w*Z�c��v���]��W5#쑻c�o�F�H��6�0��qx��+�p�_7^���;�$,���v�~�� �z=�4߯\�A��G�F�faލ�m<��|C�y�d��+:UQ���q�7���/��J��N���n�8	�	��bu�6��ь����]sJ��>���2�!3P�����h�i3ώmb�/W������+U4���Ԣ��A�s!hǔ�!٤������x}U��V��>\�)�-#�0E�B��<	�)f_�=WZ�)i�먿�Ъ-dp���*s�������b7�%M
�� �U>y����EF�G�Ė�:p�X^�}>[+Us���B.�'2@�	}�նdsLDɂ�~�k�C}��?ȕ=V�����T�n���6��K�oYN�f*�_�E0�����XE��Rze�x�xٶ@�p���ϒk�7��x�^8ָ�����}ow�r��U���P7俇c�nz[�1O�m�L��r&8h�uQ���+x�����D�o�C�����&_��8p��R�0?[ֱ|�S��0��4�,vtFoɎ�ƕ�H�����џPA@�#Y��P��"�<s�ϔ�*�� Y?���/�<��
��{o'Ô�؅h^�����\=�?'���K�WY�Hס�^H�t>��݋U� j� #������?����s�86��t���(�������w��@���aE�6�U��^uH��/���N1�4ύ7&zM�ZʦŘ���/2���*-k��MOJf��i��%(�96'����Л�����I��jT ���1~fh�-�����A�yS�!�&{N�x��B��%��s��0��涽@�j�94�l���ƛ˚H����6���mA���L�F���7\����/r/g��rO�0N(�u�Cu�o�@F�KO)Uaw�C�QgT�"fP9y^η�ۨ:�p�v�����f�o���]�v,凟�jQ�0Y_��F����چ$.H,X��M'� �6���\�X���)�LZc<�ü��0���^k��\7W_�6�j{u�~�VW%�ت����fJ�K�OC�k/�l��q�5AM�o�i*[�NibS�(۵m�����KO;��鉢�m�'2e�}&@n,Y��ߊT�]-9���(3�K ��Jvc3.��m��>X|C�{��i�Lȱ��L�w���ם�?���]i���~��5�S �&��|&��Da�R9���P��S+���ܖn;�xs3UәO'�t�,�#zV���ܮ�j�z]7�$FF���#�׉�v��!|D�g(?�ǲJtt�}��1f�z��£����l���q��b��i����$�����<�}D4+1���%t�A	��&]Нٟ�:��KE��h�D����N�w���!�)��9�0R�bH?��ð����]�G��vGވ;�G��}��ٷ��o3��_�X��jZ>u�]��L뒳�^=��|������3��:ɡ6��W&uwr���}��U�'��ڬhi[��P���#+r�(�Z���S~E��W��E��6L�:P�9��ZfS�nt5)��FD5�� #ڴ�.��_�	�#��\TKQ��*5���1�k�1��%�3s��tu���y�D,"6��5,4#��^:T�9�W�cL�y�D/5�ڤ���1t�WL�4���FA��?QN��V�`��w�+tEh!��a��VC����5�����%G$�f��.���̤�W�l�U��Y�G��?��S�gH��d��I��'_��LĲ��`r��9T��!υ�b���e��̶�e��p�m�I-�G�}�����vE"#K������.�.��J-3(�,^���cH��,�Ob�< n<;y	~��3�<�w��X~]1�F_����4�X�9����v\=��ԩt�=a1.�n�eS�-������_�BQ��\]��/��X��#<�Dh�;�3/���&���Q���ɫ�C�zsb��mД�� Ьҁ�� wt�$��8���q��r�>��4���dg#�|�e�����Qqe�>�k�=hK+�Z�-��].(��QI��$�Zx��G�}�&���Nҩ�vz}�ی����	�챿k櫺�I	���D���x�F�^|�;��j]�b�G�*����r�4<�\$�hj6��A�k�M؆k�G�8�rra�]�	Dq\xo��b���ft�f���O����E*��M�I&�zw�'\pۅ�->f�*�VqO����*P����jy}=w�lFbۆ(� Vs	Pр�/���ב���H)y��ȣ[��Xhу7Дj/$O��D�zZ��=(�z]�g�X�h��Q���@ϟ�jmr)���J���̭��>�앿tp�;�n�Xgd�IdX�bK5:�����Dpd��M��2aW�����'��^Ċ����:B5%�d�m�d��1b�k�2y�a]�|����FAhs�I�)/wب?U��xv�R&ݤ�'?�l��Z�B ���gڙ��c��$��n��u}.��b%���9�+Rn-�
��-p�~6v��kX	��[v�h�����g �'}�gU�^2��Dq��K���Nś��-����>���⭁�>N�}%RP4$0�ҿ���L*�Ռ=\���e�rr���Q�J�U�n":������O,���lJ�����T녬��P����W{6���d"�%ۆGSd
�-���M4�t�|��A�t��B�+n
�<O[�\H(KÜ$���H9D��JzSS3�K�d�G~I��Ю�;#a��s��U7&��Z�+ĝzm�R�����kQ�fM�n8zc��S�z�K�V>��q���$�j����Ο�D.��e,��o`P"�m��)RatT +�5U��k�������;A�dk����$�g��c� �k|㯎���B�����=u���A����.sQp�A9���P�����@���06n��]g#�|�͛��ϯ�oo�_����V�((��2��Y�}YrͶV�YK�g�o��V
��ht�9�-c���9[�Vɤ	,
��qK3ӯ�Gƿu�)�8W���L�͚�}��>*O��!�0�o[��
o�S[��ƧR����/�,_b_�~�'$���6W���#�F����r�߸;�R0�ªN'�j�(րVO�G��&��kO�@����ۅ<�b��������N��c�v.����f=g����ř����\��,E;m��!Jx�B1��sW��J��j���c>7�M����H�~�Qq�:�gr�s*a���|���X��i�˝�f"���,<�͍�|1��Z���nZ�X2$�*��yr5:۝J���}����1M�x�ۮ��u��]�Xvp)O}:��$�[���r���/z�q���AZ�~�m�6s5�ܤ��y,H�F�/�	���ᢹu�r��PPY�|N�Lv^1������_
w�ZFDڶ_H����c�I����������P����wHf�O�*��{^�h"��9d^���� GT4e�����G��_M�k��D���\k�����&�a�;NX���T�
P�;y�7��9��JMZ�.�l'��������yF5�m{��{� U�H$ҥ�#M!�!t� �*-@B�7AҥB(�TiPAA=�s߹���w������{��{�Y�k�9�|��_XZ�|Q��YJ��i�@������-�
c�d�讹�u��Z���NB��/�`[eh��ìD�����?ڳ]n�?�
���p§g�f��@9k���a�@����_�ت%3�m��i�%����r^�
�����`�x��e�����R�\�ʲ�k�TY�&F!x�MVD�Gk\e���g�d4���N�vٲ^~�Q�_x<J�.j%�i���8CĢP`Z��n���PS׳�B�z��
�uֶis5�F�����*���̓z�沅�4��|��"���?s�V��������> ��eh����|Mjn+���K�3wA�Tf0�)��8��DF�)G��iH-�/��� ���ͽѯ~���K�&�.�_�U�˸;+w��s*�>�z���JE����ͦ%����7U����ɀp3)�8��4'�D�\��OӘ��-�A��.T�2H��X��ڣ
�Bi7u�F�
�n�;��l��
	UMV���&��.�O:�%6�C�
��b�+O�`$��4���Ga�	��b�V'�G����za�n���ć�4�����z��e����3���h�����ɤ8���;�n�Y	j<:��m����ؖ�[R�SL�[�=?�]�ܮ�p��5"Zt�X,9vts�P/��vn{)&hY;.�v����xzI���O��suo2J�»g�:����c5�ێ�{��:><������S3L#6����5��F�R&r5n]��Gi=Vd9�> =Ɩ�����t�����wX�˝ԓ7:Ieh��Z��T?����{�~�N7{���u\����-�˄�w�3���7��d��ʒ��g	�2p�X#��3@���-���>�_�~:sOt�QZ����.uC�������:�J#�,��X�\�I��
�����s���}����
��P�˼�f�7"	���_r7�o�ru>z�����Ԭ4ƭ�A>S�_U�ۻ��\l'˹g��'�	���K-���o��]mN���\n���F�8�\s)��|���PZƟ�����ݗ5Ԝ��o��h���2Z�ꚇs���q�uNw~���*�A
QU���]��<F?���O�_)	�0TbC[���6ɘ���+��/Dl����3�Ub�ˮI)��pb�=����2ݾUo>$;Ս��ԫ��Y���1贙he{S�y����6SD�?��^�"J��o�"�C<�Ct�xG)�����վ6�U���2l��ِ��Ρi����hpשnI�9I̗n�������Q�9ֹx�YE%ҙ('r��ad{��|���G4��A�H����ڎ����'�q��İ �ʱ����5�c=EZ�J��m~�*X/�2���&f4=��5k$�#Ө�#�0��\���QVl��ʶ��r[{��3���ǖ���v�J��1�N˚�;�+�VFI���j{��d5
�2�tx�յr9�U�1� Cn�7t`CD�۩�BDJ�d>��r�4�`�V�94z��XfF���@q�h^F̭A����N}Lj�����O^E��f%�\��*�A�s?=7�4�ݵr��i?d���<���βJ_0��}J�ˤ������+!��7^�/g@�X���/T�-��	g��0׵����(scay~�f(Ys2��+��o�'�N�Ϯ�v����Pm�Wv���kV��P�*�=�6��`��m^�����z��煈>GgLϖ�_s޶�g�bQc���He���^��fF(4������Osʚ��-�������<J�/�Aޙ�d��[�+�C8�$��;��T8�����8�͟���
��u�iƎ�6p���0�+��x��DAIU䆂ȱ6��BG�i�V���ٖ��FdyD�oz�ds@,a4Q4�eX)���x�߄"S���^8,��?���-r�u��Q��p�8���p��ʢ����Q���WKF{�����Zk޷!����.<M��
ň n(|#����A��sDEsS㛑��4�Vx�6P\�NO��%l�礯j�K�;O���V�G)��s������.. +ֶ)��Φ+�`�3���8�7�}��CQ�G[�B����;bΓh�k��Ǉ}��Z1��ω��F�q���q�c�ue���tR'���w	9���4O��އ�r�\�@�@H>RV�8k�!tN�F>2����A����&\��]��U�Wn�r�´M{�X��#3B�n��s�
���W��Y[���îV+ҏ�Ï��WlW.�ה�z���//wf��w���-��ͅZUqɱR6��5��n�ԇ�U�q���@)ӎo�m߲S�JL"N���	�>xÒu�x�������n�빝� ի�q��C@)�\��{:���5���~�Aˌp�+6g��/6�һj8c����N�1��Q���Y+����*t'Ӧg���f�61	x��/�ɟ"i�x�덁)|(��DQ�*��e1=�CZ]=>� Z)%=Y�T�@�T�m�X�a�-!:�T%w��<C��0���[�d�uӐ��w-��-�Ĝ/ !�8գ<]��<�H�TA�,\�ա��^�0�>@yR"v��o��d8�yE�����
��0&(�H8N��x����8��݌��oD2�d��3���ɏ�Z��/�]�wE(6 �aC��f�3�WWo(j=5���GZ�p��b��vg�5S�4���2��.���h)~���RP�T<����)D8!�0G!b��Ÿ���4�XF��.��Uڇ
�K��ڮfD�<���1����k�����놇�\w1���0F�i,+J5�rß7����2�Ԗytc>�y0Zy�
T����$E�|j|-�/�x����:��<X�mS�`ȱo��ʘQ<���(SY�E�!9i0�0h}�!��"y���f�X\�����x�m����r��
پs2��n��ou&��ȬL��4{;���2+�;J��^g6�vr-�hP�,�$�;�h �8���X���O��v��Ҝ�"��4X<���b{�t�& ���7^kwGx1H�@�>�^ӧ���"�_p�g:�,=��a齣�&%SP��ald�T����H�y��Q�Gyٹ3�-�^�Q�R�bΉ�t���/k��_j���~8�Ɉ�j��p D�(��~��~�_�n�n��Q�$³�}��T�x?���	���{u/���;rq*E?9�B�~��V��u�wBUGu?/Eى�]}�TD)�y�e�D�P�ȯ���f�ʗ�8�U�o�OB�z�>UaD�EyȇH��"�R�IGL��nS�C�!|4�ҿ��[`8�x� Ѷ��,����ª^mi�erT��F�?\�g����A��`�x6|�s���u��!a��,I�"}0�{�K�N���G���Γ�:���%~)4|}�f}�Ž�;{���L�a	k�R�RB�����0���lo�>1�$"�k��=���B�7�)������i��w �7; W#"ц�x�)�$��D5dUS��� �<��(T���� I�#%� 'X��X/0�q���WL^���Z��+hM5��1�ź;���1a9��S��E�;tm|���S��6`�WO]�sY &�52���r�8g_�M���GvŅ�˂o'�A�;Z|4�e`"��L�A+GD�M#\���R`�NE# W�l���I.�z�s7�}���;w���u9<�e�� k�{��j5�&��,X4g~�J[*�~,��0Y���4��D�>l���f��
�h���M�Fւ,v9m���Y�;�կt�h;/GZё6�ɋ+$����L��2��6��=�P�t�>wp�ېu[GZ��7�i���޵�(��oi��D�!��	�yX�9A���d^��<�\gfv��&���j��8G6�M-'k�����,9��7!��nB�iS3�E�i^�1�Әi4�
�%;Ʌ��&�yA�9��A�����F����S�g<�!D@7CUz��#4�^[16�"Myw) zI�~��<?O�b	�4h�nDL��C�_'��g����Kme���܌�~�W�+�u�}�v�q*qC�"m��ۼLi";Ͻ��]!PWL�����;i��   ��D��=�
�<��<b�aܟ��?Q|8�œ���9=��i-� ��ȝ�叨�<<S��r��%�/i��66|�&��M�t�7�����?�o�w�Ż#�_%��Y��F�*�W��&$n�9���N��ԃ h����`�����윱k� ��:9<�+p��� q�R�98����őzn�M��~�+�僙ÃF�PMR�/�i2�PP���[э>�Nr7��]�7�U�z���0�ބ�d�{��˩FA��>��y=ߢ�a���Ұj��&�wYa7M�xG@hʒ�G��WT!��za��W�����q6�?��,��{�ޱ�9=�<x��r<B��]�����/��+]W!��)�)y ��;�:��R0��u�7���N�.�YϨb����u�F�l^6��m�t`����;�U�ͫ_n��w�e��\��]�fMY��.�n��j���NhC��\R�N�0J�\avu�׹����H���b��?�E�$}@X��@I�ڏ<b�ǖ~:��)o�����M[�~x ��n2H�ur�ECǽ�{�4CN"�|������R���?IJ����^�~��n�
1�����P�a�?�������v���zqC.�,r��a�e�f�2�sj�GX��a&uk��+��8���B>�� 0�>8��Jc���ǹ��h��T�o��njϙB�.ٟ�l��&���ZB�$	��I��#\�+Y����S���n/7�x�TB�����v�Ȗ`����9]�>U�N�f�{�
�	X��H�Cs�Į�{����Q��r��X.�?�o�����zz�TG�Ν	��ʞ�*˽j���F&�������GOY#�?��?e#H����'��!E���f�&�36NL��BfI=�oړ�XrR�M��>TK��C�%qcԌ\`z���lٍ�ҵ�ނ���k�I�*�����:ux�ڃOK��P��5%��a�U���,y7&�P�u�+�^�U�0���J'�O8���Fp^_`v����P(��Au�9\��`���\:}xx��8! �7f��dM�"�̰��h5�� 'o�G�#�+eg��]H�F0���'E�~���
,�Є,�&�*�`�;i���B��?'[�7�C�*��29H��B�m\zJ �^�xꑠ6�C���a6�D��+����1Y�X��/�M���M����*�TgGߞ�Hu^0ͷ�7`d�i��_���ӳF>!Ƅ������h�gp芈3����"KO �s?�7���a5��@l��!�4D�S���7?�wT`�۴[Gq���嶹�x��e��W5y^7�>4��)@��os��_���&���ݐ�3*BHaz�'��>^�l�}m��^��\]MV���(�ـaM�%=XO�ϒ�������ySKH����7*�s�Z5������0C;�g�?(<�'㛩��A�b�_�/� �_�O'5��a����:�Z�˟L��;���x7&g�Tf����Q)dܡ�$�H���<���|�^�@7,�G�;����e��\vK|�q�C�~����0=��D��|~NO{+����f���C��Gh�����D�<�`�Ps�i�dj4X��bb���0�@�B6�i�|�g���D�Q�y��;�?[ �E4�e�z ,%��6go��Wq TT��Τ�ms��@9�{��&4��'����f�x}��pڭUL� S��a��Otb���� �+=���T��2�0͠ռ��<����B�P����]5�'C��ҹ�o�#���O�k��nQ4 H��P�:�����w���қ�o��A��� PK   �fW�X3��  �     jsons/user_defined.json��]o�0��J�k@�$&wS�&4��B��)��0�'j3����>�,mV�
�%>�{�_s ;`	�Z��(�9p�oaj��@zȞ�mڧ�`��p��K��hsUkcӲ�;m�6<؞7�ߞ[��&�@`HsQ3��\��O27�H���<(
ۧ�s.]6��
BQgFV�Iދ�/2����Y�l]%U�
����P�U��W��#�{�G�۴��F?c�����ⴐV�_����<n�T�~s}��e��V�}%b���|!�<N0�6K�T�C[�LRї|]�@�\�!��g IY_���4$��F�t�n{����mO��{��ѕ0�<���H��̋������(�bEJ-|�\��ХIR���%&�3NS��a�)�'X#� �kV��͵"A�����8<��[V��9ND���_��vG�6@&����^��!�ף:@���M<�^W���-ūϣ@X���S��C����m�PK
   �fWV9!M�  A                  cirkitFile.jsonPK
   �eWK��"� I� /               images/4354f621-4db0-4aaf-904c-1fa28584b36b.jpgPK
   s�eWV(j�Y lw /             95 images/89e20355-1f0c-41de-86ac-b21eed32d9ff.jpgPK
   �fW�X3��  �               d� jsons/user_defined.jsonPK      <  z�   